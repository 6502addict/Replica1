library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity INTBASIC is
    port (
        clock:    in std_logic;
        cs_n:     in std_logic;
        address:  in std_logic_vector(12 downto 0);
        data_out: out std_logic_vector(7 downto 0)
    );
end entity;

architecture rtl of INTBASIC is
    -- ROM from $E000 to $FFFF (8192 bytes)
    type rom_type is array(0 to 8191) of std_logic_vector(7 downto 0);
    constant rom : rom_type := (
        X"4C", X"B0", X"E2", X"AD", X"11", X"D0", X"10", X"FB", 
        X"AD", X"10", X"D0", X"60", X"8A", X"29", X"20", X"F0", 
        X"23", X"A9", X"A0", X"85", X"E4", X"4C", X"C9", X"E3", 
        X"A9", X"20", X"C5", X"24", X"B0", X"0C", X"A9", X"8D", 
        X"A0", X"07", X"20", X"C9", X"E3", X"A9", X"A0", X"88", 
        X"D0", X"F8", X"A0", X"00", X"B1", X"E2", X"E6", X"E2", 
        X"D0", X"02", X"E6", X"E3", X"60", X"20", X"15", X"E7", 
        X"20", X"76", X"E5", X"A5", X"E2", X"C5", X"E6", X"A5", 
        X"E3", X"E5", X"E7", X"B0", X"EF", X"20", X"6D", X"E0", 
        X"4C", X"3B", X"E0", X"A5", X"CA", X"85", X"E2", X"A5", 
        X"CB", X"85", X"E3", X"A5", X"4C", X"85", X"E6", X"A5", 
        X"4D", X"85", X"E7", X"D0", X"DE", X"20", X"15", X"E7", 
        X"20", X"6D", X"E5", X"A5", X"E4", X"85", X"E2", X"A5", 
        X"E5", X"85", X"E3", X"B0", X"C7", X"86", X"D8", X"A9", 
        X"A0", X"85", X"FA", X"20", X"2A", X"E0", X"98", X"85", 
        X"E4", X"20", X"2A", X"E0", X"AA", X"20", X"2A", X"E0", 
        X"20", X"1B", X"E5", X"20", X"18", X"E0", X"84", X"FA", 
        X"AA", X"10", X"18", X"0A", X"10", X"E9", X"A5", X"E4", 
        X"D0", X"03", X"20", X"11", X"E0", X"8A", X"20", X"C9", 
        X"E3", X"A9", X"25", X"20", X"1A", X"E0", X"AA", X"30", 
        X"F5", X"85", X"E4", X"C9", X"01", X"D0", X"05", X"A6", 
        X"D8", X"4C", X"CD", X"E3", X"48", X"84", X"CE", X"A2", 
        X"ED", X"86", X"CF", X"C9", X"51", X"90", X"04", X"C6", 
        X"CF", X"E9", X"50", X"48", X"B1", X"CE", X"AA", X"88", 
        X"B1", X"CE", X"10", X"FA", X"E0", X"C0", X"B0", X"04", 
        X"E0", X"00", X"30", X"F2", X"AA", X"68", X"E9", X"01", 
        X"D0", X"E9", X"24", X"E4", X"30", X"03", X"20", X"F8", 
        X"EF", X"B1", X"CE", X"10", X"10", X"AA", X"29", X"3F", 
        X"85", X"E4", X"18", X"69", X"A0", X"20", X"C9", X"E3", 
        X"88", X"E0", X"C0", X"90", X"EC", X"20", X"0C", X"E0", 
        X"68", X"C9", X"5D", X"F0", X"A4", X"C9", X"28", X"D0", 
        X"8A", X"F0", X"9E", X"20", X"18", X"E1", X"95", X"50", 
        X"D5", X"78", X"90", X"11", X"A0", X"2B", X"4C", X"E0", 
        X"E3", X"20", X"34", X"EE", X"D5", X"50", X"90", X"F4", 
        X"20", X"E4", X"EF", X"95", X"78", X"4C", X"23", X"E8", 
        X"20", X"34", X"EE", X"F0", X"E7", X"38", X"E9", X"01", 
        X"60", X"20", X"18", X"E1", X"95", X"50", X"18", X"F5", 
        X"78", X"4C", X"02", X"E1", X"A0", X"14", X"D0", X"D6", 
        X"20", X"18", X"E1", X"E8", X"B5", X"50", X"85", X"DA", 
        X"65", X"CE", X"48", X"A8", X"B5", X"78", X"85", X"DB", 
        X"65", X"CF", X"48", X"C4", X"CA", X"E5", X"CB", X"B0", 
        X"E3", X"A5", X"DA", X"69", X"FE", X"85", X"DA", X"A9", 
        X"FF", X"A8", X"65", X"DB", X"85", X"DB", X"C8", X"B1", 
        X"DA", X"D9", X"CC", X"00", X"D0", X"0F", X"98", X"F0", 
        X"F5", X"68", X"91", X"DA", X"99", X"CC", X"00", X"88", 
        X"10", X"F7", X"E8", X"60", X"EA", X"A0", X"80", X"D0", 
        X"95", X"A9", X"00", X"20", X"0A", X"E7", X"A0", X"02", 
        X"94", X"78", X"20", X"0A", X"E7", X"A9", X"BF", X"20", 
        X"C9", X"E3", X"A0", X"00", X"20", X"9E", X"E2", X"94", 
        X"78", X"EA", X"EA", X"EA", X"B5", X"51", X"85", X"CE", 
        X"B5", X"79", X"85", X"CF", X"E8", X"E8", X"20", X"BC", 
        X"E1", X"B5", X"4E", X"D5", X"76", X"B0", X"15", X"F6", 
        X"4E", X"A8", X"B1", X"CE", X"B4", X"50", X"C4", X"E4", 
        X"90", X"04", X"A0", X"83", X"D0", X"C1", X"91", X"DA", 
        X"F6", X"50", X"90", X"E5", X"B4", X"50", X"8A", X"91", 
        X"DA", X"E8", X"E8", X"60", X"B5", X"51", X"85", X"DA", 
        X"38", X"E9", X"02", X"85", X"E4", X"B5", X"79", X"85", 
        X"DB", X"E9", X"00", X"85", X"E5", X"A0", X"00", X"B1", 
        X"E4", X"18", X"E5", X"DA", X"85", X"E4", X"60", X"B5", 
        X"53", X"85", X"CE", X"B5", X"7B", X"85", X"CF", X"B5", 
        X"51", X"85", X"DA", X"B5", X"79", X"85", X"DB", X"E8", 
        X"E8", X"E8", X"A0", X"00", X"94", X"78", X"94", X"A0", 
        X"C8", X"94", X"50", X"B5", X"4D", X"D5", X"75", X"08", 
        X"48", X"B5", X"4F", X"D5", X"77", X"90", X"07", X"68", 
        X"28", X"B0", X"02", X"56", X"50", X"60", X"A8", X"B1", 
        X"CE", X"85", X"E4", X"68", X"A8", X"28", X"B0", X"F3", 
        X"B1", X"DA", X"C5", X"E4", X"D0", X"ED", X"F6", X"4F", 
        X"F6", X"4D", X"B0", X"D7", X"20", X"D7", X"E1", X"4C", 
        X"36", X"E7", X"20", X"54", X"E2", X"06", X"CE", X"26", 
        X"CF", X"90", X"0D", X"18", X"A5", X"E6", X"65", X"DA", 
        X"85", X"E6", X"A5", X"E7", X"65", X"DB", X"85", X"E7", 
        X"88", X"F0", X"09", X"06", X"E6", X"26", X"E7", X"10", 
        X"E4", X"4C", X"7E", X"E7", X"A5", X"E6", X"20", X"08", 
        X"E7", X"A5", X"E7", X"95", X"A0", X"06", X"E5", X"90", 
        X"28", X"4C", X"6F", X"E7", X"A9", X"55", X"85", X"E5", 
        X"20", X"5B", X"E2", X"A5", X"CE", X"85", X"DA", X"A5", 
        X"CF", X"85", X"DB", X"20", X"15", X"E7", X"84", X"E6", 
        X"84", X"E7", X"A5", X"CF", X"10", X"09", X"CA", X"06", 
        X"E5", X"20", X"6F", X"E7", X"20", X"15", X"E7", X"A0", 
        X"10", X"60", X"20", X"6C", X"EE", X"F0", X"C5", X"FF", 
        X"C9", X"84", X"D0", X"02", X"46", X"F8", X"C9", X"DF", 
        X"F0", X"11", X"C9", X"9B", X"F0", X"06", X"99", X"00", 
        X"02", X"C8", X"10", X"0A", X"A0", X"8B", X"20", X"C4", 
        X"E3", X"A0", X"01", X"88", X"30", X"F6", X"20", X"03", 
        X"E0", X"EA", X"EA", X"20", X"C9", X"E3", X"C9", X"8D", 
        X"D0", X"D6", X"A9", X"DF", X"99", X"00", X"02", X"60", 
        X"20", X"D3", X"EF", X"20", X"CD", X"E3", X"46", X"D9", 
        X"A9", X"BE", X"20", X"C9", X"E3", X"A0", X"00", X"84", 
        X"FA", X"24", X"F8", X"10", X"0C", X"A6", X"F6", X"A5", 
        X"F7", X"20", X"1B", X"E5", X"A9", X"A0", X"20", X"C9", 
        X"E3", X"A2", X"FF", X"9A", X"20", X"9E", X"E2", X"84", 
        X"F1", X"8A", X"85", X"C8", X"A2", X"20", X"20", X"91", 
        X"E4", X"A5", X"C8", X"69", X"00", X"85", X"E0", X"A9", 
        X"00", X"AA", X"69", X"02", X"85", X"E1", X"A1", X"E0", 
        X"29", X"F0", X"C9", X"B0", X"F0", X"03", X"4C", X"83", 
        X"E8", X"A0", X"02", X"B1", X"E0", X"99", X"CD", X"00", 
        X"88", X"D0", X"F8", X"20", X"8A", X"E3", X"A5", X"F1", 
        X"E5", X"C8", X"C9", X"04", X"F0", X"A8", X"91", X"E0", 
        X"A5", X"CA", X"F1", X"E0", X"85", X"E4", X"A5", X"CB", 
        X"E9", X"00", X"85", X"E5", X"A5", X"E4", X"C5", X"CC", 
        X"A5", X"E5", X"E5", X"CD", X"90", X"45", X"A5", X"CA", 
        X"F1", X"E0", X"85", X"E6", X"A5", X"CB", X"E9", X"00", 
        X"85", X"E7", X"B1", X"CA", X"91", X"E6", X"E6", X"CA", 
        X"D0", X"02", X"E6", X"CB", X"A5", X"E2", X"C5", X"CA", 
        X"A5", X"E3", X"E5", X"CB", X"B0", X"E0", X"B5", X"E4", 
        X"95", X"CA", X"CA", X"10", X"F9", X"B1", X"E0", X"A8", 
        X"88", X"B1", X"E0", X"91", X"E6", X"98", X"D0", X"F8", 
        X"24", X"F8", X"10", X"09", X"B5", X"F7", X"75", X"F5", 
        X"95", X"F7", X"E8", X"F0", X"F7", X"10", X"7E", X"00", 
        X"00", X"00", X"00", X"A0", X"14", X"D0", X"71", X"20", 
        X"15", X"E7", X"A5", X"E2", X"85", X"E6", X"A5", X"E3", 
        X"85", X"E7", X"20", X"75", X"E5", X"A5", X"E2", X"85", 
        X"E4", X"A5", X"E3", X"85", X"E5", X"D0", X"0E", X"20", 
        X"15", X"E7", X"20", X"6D", X"E5", X"A5", X"E6", X"85", 
        X"E2", X"A5", X"E7", X"85", X"E3", X"A0", X"00", X"A5", 
        X"CA", X"C5", X"E4", X"A5", X"CB", X"E5", X"E5", X"B0", 
        X"16", X"A5", X"E4", X"D0", X"02", X"C6", X"E5", X"C6", 
        X"E4", X"A5", X"E6", X"D0", X"02", X"C6", X"E7", X"C6", 
        X"E6", X"B1", X"E4", X"91", X"E6", X"90", X"E0", X"A5", 
        X"E6", X"85", X"CA", X"A5", X"E7", X"85", X"CB", X"60", 
        X"20", X"C9", X"E3", X"C8", X"B9", X"00", X"EB", X"30", 
        X"F7", X"C9", X"8D", X"D0", X"06", X"A9", X"00", X"85", 
        X"24", X"A9", X"8D", X"E6", X"24", X"2C", X"12", X"D0", 
        X"30", X"FB", X"8D", X"12", X"D0", X"60", X"A0", X"06", 
        X"20", X"D3", X"EE", X"24", X"D9", X"30", X"03", X"4C", 
        X"B6", X"E2", X"4C", X"9A", X"EB", X"2A", X"69", X"A0", 
        X"DD", X"00", X"02", X"D0", X"53", X"B1", X"FE", X"0A", 
        X"30", X"06", X"88", X"B1", X"FE", X"30", X"29", X"C8", 
        X"86", X"C8", X"98", X"48", X"A2", X"00", X"A1", X"FE", 
        X"AA", X"4A", X"49", X"48", X"11", X"FE", X"C9", X"C0", 
        X"90", X"01", X"E8", X"C8", X"D0", X"F3", X"68", X"A8", 
        X"8A", X"4C", X"C0", X"E4", X"E6", X"F1", X"A6", X"F1", 
        X"F0", X"BC", X"9D", X"00", X"02", X"60", X"A6", X"C8", 
        X"A9", X"A0", X"E8", X"DD", X"00", X"02", X"B0", X"FA", 
        X"B1", X"FE", X"29", X"3F", X"4A", X"D0", X"B6", X"BD", 
        X"00", X"02", X"B0", X"06", X"69", X"3F", X"C9", X"1A", 
        X"90", X"6F", X"69", X"4F", X"C9", X"0A", X"90", X"69", 
        X"A6", X"FD", X"C8", X"B1", X"FE", X"29", X"E0", X"C9", 
        X"20", X"F0", X"7A", X"B5", X"A8", X"85", X"C8", X"B5", 
        X"D1", X"85", X"F1", X"88", X"B1", X"FE", X"0A", X"10", 
        X"FA", X"88", X"B0", X"38", X"0A", X"30", X"35", X"B4", 
        X"58", X"84", X"FF", X"B4", X"80", X"E8", X"10", X"DA", 
        X"F0", X"B3", X"C9", X"7E", X"B0", X"22", X"CA", X"10", 
        X"04", X"A0", X"06", X"10", X"29", X"94", X"80", X"A4", 
        X"FF", X"94", X"58", X"A4", X"C8", X"94", X"A8", X"A4", 
        X"F1", X"94", X"D1", X"29", X"1F", X"A8", X"B9", X"20", 
        X"EC", X"0A", X"A8", X"A9", X"76", X"2A", X"85", X"FF", 
        X"D0", X"01", X"C8", X"C8", X"86", X"FD", X"B1", X"FE", 
        X"30", X"84", X"D0", X"05", X"A0", X"0E", X"4C", X"E0", 
        X"E3", X"C9", X"03", X"B0", X"C3", X"4A", X"A6", X"C8", 
        X"E8", X"BD", X"00", X"02", X"90", X"04", X"C9", X"A2", 
        X"F0", X"0A", X"C9", X"DF", X"F0", X"06", X"86", X"C8", 
        X"20", X"1C", X"E4", X"C8", X"88", X"A6", X"FD", X"B1", 
        X"FE", X"88", X"0A", X"10", X"CF", X"B4", X"58", X"84", 
        X"FF", X"B4", X"80", X"E8", X"B1", X"FE", X"29", X"9F", 
        X"D0", X"ED", X"85", X"F2", X"85", X"F3", X"98", X"48", 
        X"86", X"FD", X"B4", X"D0", X"84", X"C9", X"18", X"A9", 
        X"0A", X"85", X"F9", X"A2", X"00", X"C8", X"B9", X"00", 
        X"02", X"29", X"0F", X"65", X"F2", X"48", X"8A", X"65", 
        X"F3", X"30", X"1C", X"AA", X"68", X"C6", X"F9", X"D0", 
        X"F2", X"85", X"F2", X"86", X"F3", X"C4", X"F1", X"D0", 
        X"DE", X"A4", X"C9", X"C8", X"84", X"F1", X"20", X"1C", 
        X"E4", X"68", X"A8", X"A5", X"F3", X"B0", X"A9", X"A0", 
        X"00", X"10", X"8B", X"85", X"F3", X"86", X"F2", X"A2", 
        X"04", X"86", X"C9", X"A9", X"B0", X"85", X"F9", X"A5", 
        X"F2", X"DD", X"63", X"E5", X"A5", X"F3", X"FD", X"68", 
        X"E5", X"90", X"0D", X"85", X"F3", X"A5", X"F2", X"FD", 
        X"63", X"E5", X"85", X"F2", X"E6", X"F9", X"D0", X"E7", 
        X"A5", X"F9", X"E8", X"CA", X"F0", X"0E", X"C9", X"B0", 
        X"F0", X"02", X"85", X"C9", X"24", X"C9", X"30", X"04", 
        X"A5", X"FA", X"F0", X"0B", X"20", X"C9", X"E3", X"24", 
        X"F8", X"10", X"04", X"99", X"00", X"02", X"C8", X"CA", 
        X"10", X"C1", X"60", X"01", X"0A", X"64", X"E8", X"10", 
        X"00", X"00", X"00", X"03", X"27", X"A5", X"CA", X"85", 
        X"E6", X"A5", X"CB", X"85", X"E7", X"E8", X"A5", X"E7", 
        X"85", X"E5", X"A5", X"E6", X"85", X"E4", X"C5", X"4C", 
        X"A5", X"E5", X"E5", X"4D", X"B0", X"26", X"A0", X"01", 
        X"B1", X"E4", X"E5", X"CE", X"C8", X"B1", X"E4", X"E5", 
        X"CF", X"B0", X"19", X"A0", X"00", X"A5", X"E6", X"71", 
        X"E4", X"85", X"E6", X"90", X"03", X"E6", X"E7", X"18", 
        X"C8", X"A5", X"CE", X"F1", X"E4", X"C8", X"A5", X"CF", 
        X"F1", X"E4", X"B0", X"CA", X"60", X"46", X"F8", X"A5", 
        X"4C", X"85", X"CA", X"A5", X"4D", X"85", X"CB", X"A5", 
        X"4A", X"85", X"CC", X"A5", X"4B", X"85", X"CD", X"A9", 
        X"00", X"85", X"FB", X"85", X"FC", X"85", X"FE", X"A9", 
        X"00", X"85", X"1D", X"60", X"A5", X"D0", X"69", X"05", 
        X"85", X"D2", X"A5", X"D1", X"69", X"00", X"85", X"D3", 
        X"A5", X"D2", X"C5", X"CA", X"A5", X"D3", X"E5", X"CB", 
        X"90", X"03", X"4C", X"6B", X"E3", X"A5", X"CE", X"91", 
        X"D0", X"A5", X"CF", X"C8", X"91", X"D0", X"A5", X"D2", 
        X"C8", X"91", X"D0", X"A5", X"D3", X"C8", X"91", X"D0", 
        X"A9", X"00", X"C8", X"91", X"D0", X"C8", X"91", X"D0", 
        X"A5", X"D2", X"85", X"CC", X"A5", X"D3", X"85", X"CD", 
        X"A5", X"D0", X"90", X"43", X"85", X"CE", X"84", X"CF", 
        X"20", X"FF", X"E6", X"30", X"0E", X"C9", X"40", X"F0", 
        X"0A", X"4C", X"28", X"E6", X"06", X"C9", X"49", X"D0", 
        X"07", X"A9", X"49", X"85", X"CF", X"20", X"FF", X"E6", 
        X"A5", X"4B", X"85", X"D1", X"A5", X"4A", X"85", X"D0", 
        X"C5", X"CC", X"A5", X"D1", X"E5", X"CD", X"B0", X"94", 
        X"B1", X"D0", X"C8", X"C5", X"CE", X"D0", X"06", X"B1", 
        X"D0", X"C5", X"CF", X"F0", X"0E", X"C8", X"B1", X"D0", 
        X"48", X"C8", X"B1", X"D0", X"85", X"D1", X"68", X"A0", 
        X"00", X"F0", X"DB", X"A5", X"D0", X"69", X"03", X"20", 
        X"0A", X"E7", X"A5", X"D1", X"69", X"00", X"95", X"78", 
        X"A5", X"CF", X"C9", X"40", X"D0", X"1C", X"88", X"98", 
        X"20", X"0A", X"E7", X"88", X"94", X"78", X"A0", X"03", 
        X"F6", X"78", X"C8", X"B1", X"D0", X"30", X"F9", X"10", 
        X"09", X"A9", X"00", X"85", X"D4", X"85", X"D5", X"A2", 
        X"20", X"48", X"A0", X"00", X"B1", X"E0", X"10", X"18", 
        X"0A", X"30", X"81", X"20", X"FF", X"E6", X"20", X"08", 
        X"E7", X"20", X"FF", X"E6", X"95", X"A0", X"24", X"D4", 
        X"10", X"01", X"CA", X"20", X"FF", X"E6", X"B0", X"E6", 
        X"C9", X"28", X"D0", X"1F", X"A5", X"E0", X"20", X"0A", 
        X"E7", X"A5", X"E1", X"95", X"78", X"24", X"D4", X"30", 
        X"0B", X"A9", X"01", X"20", X"0A", X"E7", X"A9", X"00", 
        X"95", X"78", X"F6", X"78", X"20", X"FF", X"E6", X"30", 
        X"F9", X"B0", X"D3", X"24", X"D4", X"10", X"06", X"C9", 
        X"04", X"B0", X"D0", X"46", X"D4", X"A8", X"85", X"D6", 
        X"B9", X"98", X"E9", X"29", X"55", X"0A", X"85", X"D7", 
        X"68", X"A8", X"B9", X"98", X"E9", X"29", X"AA", X"C5", 
        X"D7", X"B0", X"09", X"98", X"48", X"20", X"FF", X"E6", 
        X"A5", X"D6", X"90", X"95", X"B9", X"10", X"EA", X"85", 
        X"CE", X"B9", X"88", X"EA", X"85", X"CF", X"20", X"FC", 
        X"E6", X"4C", X"D8", X"E6", X"6C", X"CE", X"00", X"E6", 
        X"E0", X"D0", X"02", X"E6", X"E1", X"B1", X"E0", X"60", 
        X"94", X"77", X"CA", X"30", X"03", X"95", X"50", X"60", 
        X"A0", X"66", X"4C", X"E0", X"E3", X"A0", X"00", X"B5", 
        X"50", X"85", X"CE", X"B5", X"A0", X"85", X"CF", X"B5", 
        X"78", X"F0", X"0E", X"85", X"CF", X"B1", X"CE", X"48", 
        X"C8", X"B1", X"CE", X"85", X"CF", X"68", X"85", X"CE", 
        X"88", X"E8", X"60", X"20", X"4A", X"E7", X"20", X"15", 
        X"E7", X"98", X"20", X"08", X"E7", X"95", X"A0", X"C5", 
        X"CE", X"D0", X"06", X"C5", X"CF", X"D0", X"02", X"F6", 
        X"50", X"60", X"20", X"82", X"E7", X"20", X"59", X"E7", 
        X"20", X"15", X"E7", X"24", X"CF", X"30", X"1B", X"CA", 
        X"60", X"20", X"15", X"E7", X"A5", X"CF", X"D0", X"04", 
        X"A5", X"CE", X"F0", X"F3", X"A9", X"FF", X"20", X"08", 
        X"E7", X"95", X"A0", X"24", X"CF", X"30", X"E9", X"20", 
        X"15", X"E7", X"98", X"38", X"E5", X"CE", X"20", X"08", 
        X"E7", X"98", X"E5", X"CF", X"50", X"23", X"A0", X"00", 
        X"10", X"90", X"20", X"6F", X"E7", X"20", X"15", X"E7", 
        X"A5", X"CE", X"85", X"DA", X"A5", X"CF", X"85", X"DB", 
        X"20", X"15", X"E7", X"18", X"A5", X"CE", X"65", X"DA", 
        X"20", X"08", X"E7", X"A5", X"CF", X"65", X"DB", X"70", 
        X"DD", X"95", X"A0", X"60", X"20", X"15", X"E7", X"A4", 
        X"CE", X"F0", X"05", X"88", X"A5", X"CF", X"F0", X"0C", 
        X"60", X"A5", X"24", X"09", X"07", X"A8", X"C8", X"A9", 
        X"A0", X"20", X"C9", X"E3", X"C4", X"24", X"B0", X"F7", 
        X"60", X"20", X"B1", X"E7", X"20", X"15", X"E7", X"A5", 
        X"CF", X"10", X"0A", X"A9", X"AD", X"20", X"C9", X"E3", 
        X"20", X"72", X"E7", X"50", X"EF", X"88", X"84", X"D5", 
        X"86", X"CF", X"A6", X"CE", X"20", X"1B", X"E5", X"A6", 
        X"CF", X"60", X"20", X"15", X"E7", X"A5", X"CE", X"85", 
        X"F6", X"A5", X"CF", X"85", X"F7", X"88", X"84", X"F8", 
        X"C8", X"A9", X"0A", X"85", X"F4", X"84", X"F5", X"60", 
        X"20", X"15", X"E7", X"A5", X"CE", X"A4", X"CF", X"10", 
        X"F2", X"20", X"15", X"E7", X"B5", X"50", X"85", X"DA", 
        X"B5", X"78", X"85", X"DB", X"A5", X"CE", X"91", X"DA", 
        X"C8", X"A5", X"CF", X"91", X"DA", X"E8", X"60", X"68", 
        X"68", X"24", X"D5", X"10", X"05", X"20", X"CD", X"E3", 
        X"46", X"D5", X"60", X"A0", X"FF", X"84", X"D7", X"60", 
        X"20", X"CD", X"EF", X"F0", X"07", X"A9", X"25", X"85", 
        X"D6", X"88", X"84", X"D4", X"E8", X"60", X"A5", X"CA", 
        X"A4", X"CB", X"D0", X"5A", X"A0", X"41", X"A5", X"FC", 
        X"C9", X"08", X"B0", X"5E", X"A8", X"E6", X"FC", X"A5", 
        X"E0", X"99", X"00", X"01", X"A5", X"E1", X"99", X"08", 
        X"01", X"A5", X"DC", X"99", X"10", X"01", X"A5", X"DD", 
        X"99", X"18", X"01", X"20", X"15", X"E7", X"20", X"6D", 
        X"E5", X"90", X"04", X"A0", X"37", X"D0", X"3B", X"A5", 
        X"E4", X"A4", X"E5", X"85", X"DC", X"84", X"DD", X"2C", 
        X"11", X"D0", X"30", X"4F", X"18", X"69", X"03", X"90", 
        X"01", X"C8", X"A2", X"FF", X"86", X"D9", X"9A", X"85", 
        X"E0", X"84", X"E1", X"20", X"79", X"E6", X"24", X"D9", 
        X"10", X"49", X"18", X"A0", X"00", X"A5", X"DC", X"71", 
        X"DC", X"A4", X"DD", X"90", X"01", X"C8", X"C5", X"4C", 
        X"D0", X"D1", X"C4", X"4D", X"D0", X"CD", X"A0", X"34", 
        X"46", X"D9", X"4C", X"E0", X"E3", X"A0", X"4A", X"A5", 
        X"FC", X"F0", X"F7", X"C6", X"FC", X"A8", X"B9", X"0F", 
        X"01", X"85", X"DC", X"B9", X"17", X"01", X"85", X"DD", 
        X"BE", X"FF", X"00", X"B9", X"07", X"01", X"A8", X"8A", 
        X"4C", X"7A", X"E8", X"A0", X"63", X"20", X"C4", X"E3", 
        X"A0", X"01", X"B1", X"DC", X"AA", X"C8", X"B1", X"DC", 
        X"20", X"1B", X"E5", X"4C", X"B3", X"E2", X"C6", X"FB", 
        X"A0", X"5B", X"A5", X"FB", X"F0", X"C4", X"A8", X"B5", 
        X"50", X"D9", X"1F", X"01", X"D0", X"F0", X"B5", X"78", 
        X"D9", X"27", X"01", X"D0", X"E9", X"B9", X"2F", X"01", 
        X"85", X"DA", X"B9", X"37", X"01", X"85", X"DB", X"20", 
        X"15", X"E7", X"CA", X"20", X"93", X"E7", X"20", X"01", 
        X"E8", X"CA", X"A4", X"FB", X"B9", X"67", X"01", X"95", 
        X"9F", X"B9", X"5F", X"01", X"A0", X"00", X"20", X"08", 
        X"E7", X"20", X"82", X"E7", X"20", X"59", X"E7", X"20", 
        X"15", X"E7", X"A4", X"FB", X"A5", X"CE", X"F0", X"05", 
        X"59", X"37", X"01", X"10", X"12", X"B9", X"3F", X"01", 
        X"85", X"DC", X"B9", X"47", X"01", X"85", X"DD", X"BE", 
        X"4F", X"01", X"B9", X"57", X"01", X"D0", X"87", X"C6", 
        X"FB", X"60", X"A0", X"54", X"A5", X"FB", X"C9", X"08", 
        X"F0", X"9A", X"E6", X"FB", X"A8", X"B5", X"50", X"99", 
        X"20", X"01", X"B5", X"78", X"99", X"28", X"01", X"60", 
        X"20", X"15", X"E7", X"A4", X"FB", X"A5", X"CE", X"99", 
        X"5F", X"01", X"A5", X"CF", X"99", X"67", X"01", X"A9", 
        X"01", X"99", X"2F", X"01", X"A9", X"00", X"99", X"37", 
        X"01", X"A5", X"DC", X"99", X"3F", X"01", X"A5", X"DD", 
        X"99", X"47", X"01", X"A5", X"E0", X"99", X"4F", X"01", 
        X"A5", X"E1", X"99", X"57", X"01", X"60", X"20", X"15", 
        X"E7", X"A4", X"FB", X"A5", X"CE", X"99", X"2F", X"01", 
        X"A5", X"CF", X"4C", X"66", X"E9", X"00", X"00", X"00", 
        X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
        X"00", X"00", X"00", X"AB", X"03", X"03", X"03", X"03", 
        X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", 
        X"03", X"03", X"3F", X"3F", X"C0", X"C0", X"3C", X"3C", 
        X"3C", X"3C", X"3C", X"3C", X"3C", X"30", X"0F", X"C0", 
        X"CC", X"FF", X"55", X"00", X"AB", X"AB", X"03", X"03", 
        X"FF", X"FF", X"55", X"FF", X"FF", X"55", X"CF", X"CF", 
        X"CF", X"CF", X"CF", X"FF", X"55", X"C3", X"C3", X"C3", 
        X"55", X"F0", X"F0", X"CF", X"56", X"56", X"56", X"55", 
        X"FF", X"FF", X"55", X"03", X"03", X"03", X"03", X"03", 
        X"03", X"03", X"FF", X"FF", X"FF", X"03", X"03", X"03", 
        X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", 
        X"03", X"03", X"03", X"03", X"03", X"00", X"AB", X"03", 
        X"57", X"03", X"03", X"03", X"03", X"07", X"03", X"03", 
        X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", 
        X"03", X"03", X"AA", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"17", X"FF", X"FF", X"19", X"5D", X"35", X"4B", X"F2", 
        X"EC", X"87", X"6F", X"AD", X"B7", X"E2", X"F8", X"54", 
        X"80", X"96", X"85", X"82", X"22", X"10", X"33", X"4A", 
        X"13", X"06", X"0B", X"4A", X"01", X"40", X"47", X"7A", 
        X"00", X"FF", X"23", X"09", X"5B", X"16", X"B6", X"CB", 
        X"FF", X"FF", X"FB", X"FF", X"FF", X"24", X"F6", X"4E", 
        X"59", X"50", X"00", X"FF", X"23", X"A3", X"6F", X"36", 
        X"23", X"D7", X"1C", X"22", X"C2", X"AE", X"BA", X"23", 
        X"FF", X"FF", X"21", X"30", X"1E", X"03", X"C4", X"20", 
        X"00", X"C1", X"FF", X"FF", X"FF", X"A0", X"30", X"1E", 
        X"A4", X"D3", X"B6", X"BC", X"AA", X"3A", X"01", X"50", 
        X"7E", X"D8", X"D8", X"A5", X"3C", X"FF", X"16", X"5B", 
        X"28", X"03", X"C4", X"1D", X"00", X"0C", X"4E", X"00", 
        X"3E", X"00", X"A6", X"B0", X"00", X"BC", X"C6", X"57", 
        X"8C", X"01", X"27", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"E8", X"FF", X"FF", X"E8", X"E0", X"E0", X"E0", X"EF", 
        X"EF", X"E3", X"E3", X"E5", X"E5", X"E7", X"E7", X"EE", 
        X"EF", X"EF", X"E7", X"E7", X"E2", X"EF", X"E7", X"E7", 
        X"EC", X"EC", X"EC", X"E7", X"EC", X"EC", X"EC", X"E2", 
        X"00", X"FF", X"E8", X"E1", X"E8", X"E8", X"EF", X"EB", 
        X"FF", X"FF", X"E0", X"FF", X"FF", X"EF", X"EE", X"EF", 
        X"E7", X"E7", X"00", X"FF", X"E8", X"E7", X"E7", X"E7", 
        X"E8", X"E1", X"E2", X"EE", X"EE", X"EE", X"EE", X"E8", 
        X"FF", X"FF", X"E1", X"E1", X"EF", X"EE", X"E7", X"E8", 
        X"EE", X"E7", X"FF", X"FF", X"FF", X"EE", X"E1", X"EF", 
        X"E7", X"E8", X"EF", X"EF", X"EB", X"E9", X"E8", X"E9", 
        X"E9", X"E8", X"E8", X"E8", X"E8", X"FF", X"E8", X"E8", 
        X"E8", X"EE", X"E7", X"E8", X"EF", X"EF", X"EE", X"EF", 
        X"EE", X"EF", X"EE", X"EE", X"EF", X"EE", X"EE", X"EE", 
        X"E1", X"E8", X"E8", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"BE", X"B3", X"B2", X"B7", X"B6", X"37", X"D4", X"CF", 
        X"CF", X"A0", X"CC", X"CF", X"CE", X"47", X"D3", X"D9", 
        X"CE", X"D4", X"C1", X"58", X"CD", X"C5", X"CD", X"A0", 
        X"C6", X"D5", X"CC", X"4C", X"D4", X"CF", X"CF", X"A0", 
        X"CD", X"C1", X"CE", X"D9", X"A0", X"D0", X"C1", X"D2", 
        X"C5", X"CE", X"53", X"D3", X"D4", X"D2", X"C9", X"CE", 
        X"47", X"CE", X"CF", X"A0", X"C5", X"CE", X"44", X"C2", 
        X"C1", X"C4", X"A0", X"C2", X"D2", X"C1", X"CE", X"C3", 
        X"48", X"BE", X"B8", X"A0", X"C7", X"CF", X"D3", X"D5", 
        X"C2", X"53", X"C2", X"C1", X"C4", X"A0", X"D2", X"C5", 
        X"D4", X"D5", X"D2", X"4E", X"BE", X"B8", X"A0", X"C6", 
        X"CF", X"D2", X"53", X"C2", X"C1", X"C4", X"A0", X"CE", 
        X"C5", X"D8", X"54", X"D3", X"D4", X"CF", X"D0", X"D0", 
        X"C5", X"C4", X"A0", X"C1", X"D4", X"20", X"AA", X"AA", 
        X"AA", X"20", X"A0", X"C5", X"D2", X"D2", X"0D", X"BE", 
        X"B2", X"B5", X"35", X"D2", X"C1", X"CE", X"C7", X"45", 
        X"C4", X"C9", X"4D", X"D3", X"D4", X"D2", X"A0", X"CF", 
        X"D6", X"C6", X"4C", X"DC", X"0D", X"D2", X"C5", X"D4", 
        X"D9", X"D0", X"C5", X"A0", X"CC", X"C9", X"CE", X"C5", 
        X"8D", X"3F", X"46", X"D9", X"90", X"03", X"4C", X"C3", 
        X"E8", X"A6", X"CF", X"9A", X"A6", X"CE", X"A0", X"8D", 
        X"D0", X"02", X"A0", X"99", X"20", X"C4", X"E3", X"86", 
        X"CE", X"BA", X"86", X"CF", X"A0", X"FE", X"84", X"D9", 
        X"C8", X"84", X"C8", X"20", X"99", X"E2", X"84", X"F1", 
        X"A2", X"20", X"A9", X"30", X"20", X"91", X"E4", X"E6", 
        X"D9", X"A6", X"CE", X"A4", X"C8", X"0A", X"85", X"CE", 
        X"C8", X"B9", X"00", X"02", X"C9", X"74", X"F0", X"D2", 
        X"49", X"B0", X"C9", X"0A", X"B0", X"F0", X"C8", X"C8", 
        X"84", X"C8", X"B9", X"00", X"02", X"48", X"B9", X"FF", 
        X"01", X"A0", X"00", X"20", X"08", X"E7", X"68", X"95", 
        X"A0", X"A5", X"CE", X"C9", X"C7", X"D0", X"03", X"20", 
        X"6F", X"E7", X"4C", X"01", X"E8", X"FF", X"FF", X"FF", 
        X"50", X"20", X"13", X"EC", X"D0", X"15", X"20", X"0B", 
        X"EC", X"D0", X"10", X"20", X"82", X"E7", X"20", X"6F", 
        X"E7", X"50", X"03", X"20", X"82", X"E7", X"20", X"59", 
        X"E7", X"56", X"50", X"4C", X"36", X"E7", X"FF", X"FF", 
        X"C1", X"FF", X"7F", X"D1", X"CC", X"C7", X"CF", X"CE", 
        X"C5", X"9A", X"98", X"8B", X"96", X"95", X"93", X"BF", 
        X"B2", X"32", X"2D", X"2B", X"BC", X"B0", X"AC", X"BE", 
        X"35", X"8E", X"61", X"FF", X"FF", X"FF", X"DD", X"FB", 
        X"20", X"C9", X"EF", X"15", X"4F", X"10", X"05", X"20", 
        X"C9", X"EF", X"35", X"4F", X"95", X"50", X"10", X"CB", 
        X"4C", X"C9", X"EF", X"40", X"60", X"8D", X"60", X"8B", 
        X"00", X"7E", X"8C", X"33", X"00", X"00", X"60", X"03", 
        X"BF", X"12", X"00", X"40", X"89", X"C9", X"47", X"9D", 
        X"17", X"68", X"9D", X"0A", X"00", X"40", X"60", X"8D", 
        X"60", X"8B", X"00", X"7E", X"8C", X"3C", X"00", X"00", 
        X"60", X"03", X"BF", X"1B", X"4B", X"67", X"B4", X"A1", 
        X"07", X"8C", X"07", X"AE", X"A9", X"AC", X"A8", X"67", 
        X"8C", X"07", X"B4", X"AF", X"AC", X"B0", X"67", X"9D", 
        X"B2", X"AF", X"AC", X"AF", X"A3", X"67", X"8C", X"07", 
        X"A5", X"AB", X"AF", X"B0", X"F4", X"AE", X"A9", X"B2", 
        X"B0", X"7F", X"0E", X"27", X"B4", X"AE", X"A9", X"B2", 
        X"B0", X"7F", X"0E", X"28", X"B4", X"AE", X"A9", X"B2", 
        X"B0", X"64", X"07", X"A6", X"A9", X"67", X"AF", X"B4", 
        X"AF", X"A7", X"78", X"B4", X"A5", X"AC", X"78", X"7F", 
        X"02", X"AD", X"A5", X"B2", X"67", X"A2", X"B5", X"B3", 
        X"AF", X"A7", X"EE", X"B2", X"B5", X"B4", X"A5", X"B2", 
        X"7E", X"8C", X"39", X"B4", X"B8", X"A5", X"AE", X"67", 
        X"B0", X"A5", X"B4", X"B3", X"27", X"AF", X"B4", X"07", 
        X"9D", X"19", X"B2", X"AF", X"A6", X"7F", X"05", X"37", 
        X"B4", X"B5", X"B0", X"AE", X"A9", X"7F", X"05", X"28", 
        X"B4", X"B5", X"B0", X"AE", X"A9", X"7F", X"05", X"2A", 
        X"B4", X"B5", X"B0", X"AE", X"A9", X"E4", X"AE", X"A5", 
        X"00", X"FF", X"FF", X"47", X"A2", X"A1", X"B4", X"7F", 
        X"0D", X"30", X"AD", X"A9", X"A4", X"7F", X"0D", X"23", 
        X"AD", X"A9", X"A4", X"67", X"AC", X"AC", X"A1", X"A3", 
        X"00", X"40", X"80", X"C0", X"C1", X"80", X"00", X"47", 
        X"8C", X"68", X"8C", X"DB", X"67", X"9B", X"68", X"9B", 
        X"50", X"8C", X"63", X"8C", X"7F", X"01", X"51", X"07", 
        X"88", X"29", X"84", X"80", X"C4", X"80", X"57", X"71", 
        X"07", X"88", X"14", X"ED", X"A5", X"AD", X"AF", X"AC", 
        X"ED", X"A5", X"AD", X"A9", X"A8", X"F2", X"AF", X"AC", 
        X"AF", X"A3", X"71", X"08", X"88", X"AE", X"A5", X"AC", 
        X"68", X"83", X"08", X"68", X"9D", X"08", X"71", X"07", 
        X"88", X"60", X"76", X"B4", X"AF", X"AE", X"76", X"8D", 
        X"76", X"8B", X"51", X"07", X"88", X"19", X"B8", X"A4", 
        X"AE", X"B2", X"F2", X"B3", X"B5", X"F3", X"A2", X"A1", 
        X"EE", X"A7", X"B3", X"E4", X"AE", X"B2", X"EB", X"A5", 
        X"A5", X"B0", X"51", X"07", X"88", X"39", X"81", X"C1", 
        X"4F", X"7F", X"0F", X"2F", X"00", X"51", X"06", X"88", 
        X"29", X"C2", X"0C", X"82", X"57", X"8C", X"6A", X"8C", 
        X"42", X"AE", X"A5", X"A8", X"B4", X"60", X"AE", X"A5", 
        X"A8", X"B4", X"4F", X"7E", X"1E", X"35", X"8C", X"27", 
        X"51", X"07", X"88", X"09", X"8B", X"FE", X"E4", X"AF", 
        X"AD", X"F2", X"AF", X"E4", X"AE", X"A1", X"DC", X"DE", 
        X"9C", X"DD", X"9C", X"DE", X"DD", X"9E", X"C3", X"DD", 
        X"CF", X"CA", X"CD", X"CB", X"00", X"47", X"9D", X"AD", 
        X"A5", X"AD", X"AF", X"AC", X"76", X"9D", X"AD", X"A5", 
        X"AD", X"A9", X"A8", X"E6", X"A6", X"AF", X"60", X"8C", 
        X"20", X"AF", X"B4", X"B5", X"A1", X"F2", X"AC", X"A3", 
        X"F2", X"A3", X"B3", X"60", X"8C", X"20", X"AC", X"A5", 
        X"A4", X"EE", X"B5", X"B2", X"60", X"AE", X"B5", X"B2", 
        X"F4", X"B3", X"A9", X"AC", X"60", X"8C", X"20", X"B4", 
        X"B3", X"A9", X"AC", X"7A", X"7E", X"9A", X"22", X"20", 
        X"00", X"60", X"03", X"BF", X"60", X"03", X"BF", X"1F", 
        X"20", X"B1", X"E7", X"E8", X"E8", X"B5", X"4F", X"85", 
        X"DA", X"B5", X"77", X"85", X"DB", X"B4", X"4E", X"98", 
        X"D5", X"76", X"B0", X"09", X"B1", X"DA", X"20", X"C9", 
        X"E3", X"C8", X"4C", X"0F", X"EE", X"A9", X"FF", X"85", 
        X"D5", X"60", X"E8", X"A9", X"00", X"95", X"78", X"95", 
        X"A0", X"B5", X"77", X"38", X"F5", X"4F", X"95", X"50", 
        X"4C", X"23", X"E8", X"FF", X"20", X"15", X"E7", X"A5", 
        X"CF", X"D0", X"28", X"A5", X"CE", X"60", X"20", X"34", 
        X"EE", X"A4", X"C8", X"C9", X"30", X"B0", X"21", X"C0", 
        X"28", X"B0", X"1D", X"60", X"EA", X"EA", X"20", X"34", 
        X"EE", X"60", X"EA", X"8A", X"A2", X"01", X"B4", X"CE", 
        X"94", X"4C", X"B4", X"48", X"94", X"CA", X"CA", X"F0", 
        X"F5", X"AA", X"60", X"A0", X"77", X"4C", X"E0", X"E3", 
        X"A0", X"7B", X"D0", X"F9", X"20", X"54", X"E2", X"A5", 
        X"DA", X"D0", X"07", X"A5", X"DB", X"D0", X"03", X"4C", 
        X"7E", X"E7", X"06", X"CE", X"26", X"CF", X"26", X"E6", 
        X"26", X"E7", X"A5", X"E6", X"C5", X"DA", X"A5", X"E7", 
        X"E5", X"DB", X"90", X"0A", X"85", X"E7", X"A5", X"E6", 
        X"E5", X"DA", X"85", X"E6", X"E6", X"CE", X"88", X"D0", 
        X"E1", X"60", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
        X"20", X"15", X"E7", X"6C", X"CE", X"00", X"A5", X"4C", 
        X"D0", X"02", X"C6", X"4D", X"C6", X"4C", X"A5", X"48", 
        X"D0", X"02", X"C6", X"49", X"C6", X"48", X"A0", X"00", 
        X"B1", X"4C", X"91", X"48", X"A5", X"CA", X"C5", X"4C", 
        X"A5", X"CB", X"E5", X"4D", X"90", X"E0", X"4C", X"53", 
        X"EE", X"C9", X"28", X"B0", X"9B", X"A8", X"A5", X"C8", 
        X"60", X"EA", X"EA", X"98", X"AA", X"A0", X"6E", X"20", 
        X"C4", X"E3", X"8A", X"A8", X"20", X"C4", X"E3", X"A0", 
        X"72", X"4C", X"C4", X"E3", X"20", X"15", X"E7", X"06", 
        X"CE", X"26", X"CF", X"30", X"FA", X"B0", X"DC", X"D0", 
        X"04", X"C5", X"CE", X"B0", X"D6", X"60", X"20", X"15", 
        X"E7", X"B1", X"CE", X"94", X"9F", X"4C", X"08", X"E7", 
        X"20", X"34", X"EE", X"A5", X"CE", X"48", X"20", X"15", 
        X"E7", X"68", X"91", X"CE", X"60", X"FF", X"FF", X"FF", 
        X"20", X"6C", X"EE", X"A5", X"CE", X"85", X"E6", X"A5", 
        X"CF", X"85", X"E7", X"4C", X"44", X"E2", X"20", X"E4", 
        X"EE", X"4C", X"34", X"E1", X"20", X"E4", X"EE", X"B4", 
        X"78", X"B5", X"50", X"69", X"FE", X"B0", X"01", X"88", 
        X"85", X"DA", X"84", X"DB", X"18", X"65", X"CE", X"95", 
        X"50", X"98", X"65", X"CF", X"95", X"78", X"A0", X"00", 
        X"B5", X"50", X"D1", X"DA", X"C8", X"B5", X"78", X"F1", 
        X"DA", X"B0", X"80", X"4C", X"23", X"E8", X"20", X"15", 
        X"E7", X"A5", X"4E", X"20", X"08", X"E7", X"A5", X"4F", 
        X"D0", X"04", X"C5", X"4E", X"69", X"00", X"29", X"7F", 
        X"85", X"4F", X"95", X"A0", X"A0", X"11", X"A5", X"4F", 
        X"0A", X"18", X"69", X"40", X"0A", X"26", X"4E", X"26", 
        X"4F", X"88", X"D0", X"F2", X"A5", X"CE", X"20", X"08", 
        X"E7", X"A5", X"CF", X"95", X"A0", X"4C", X"7A", X"E2", 
        X"20", X"15", X"E7", X"A4", X"CE", X"C4", X"4C", X"A5", 
        X"CF", X"E5", X"4D", X"90", X"1F", X"84", X"48", X"A5", 
        X"CF", X"85", X"49", X"4C", X"B6", X"EE", X"20", X"15", 
        X"E7", X"A4", X"CE", X"C4", X"CA", X"A5", X"CF", X"E5", 
        X"CB", X"B0", X"09", X"84", X"4A", X"A5", X"CF", X"85", 
        X"4B", X"4C", X"B7", X"E5", X"4C", X"CB", X"EE", X"EA", 
        X"EA", X"EA", X"EA", X"20", X"C9", X"EF", X"20", X"71", 
        X"E1", X"4C", X"BF", X"EF", X"20", X"03", X"EE", X"A9", 
        X"FF", X"85", X"C8", X"A9", X"74", X"8D", X"00", X"02", 
        X"60", X"20", X"36", X"E7", X"E8", X"20", X"36", X"E7", 
        X"B5", X"50", X"60", X"A9", X"00", X"85", X"4A", X"85", 
        X"4C", X"A9", X"08", X"85", X"4B", X"A9", X"10", X"85", 
        X"4D", X"4C", X"AD", X"E5", X"D5", X"78", X"D0", X"01", 
        X"18", X"4C", X"02", X"E1", X"20", X"B7", X"E5", X"4C", 
        X"36", X"E8", X"20", X"B7", X"E5", X"4C", X"5B", X"E8", 
        X"E0", X"80", X"D0", X"01", X"88", X"4C", X"0C", X"E0", 
        X"A9", X"03", X"85", X"F8", X"A9", X"20", X"85", X"FF", 
        X"A9", X"7C", X"85", X"F9", X"A2", X"1B", X"BD", X"67", 
        X"FD", X"20", X"EF", X"FF", X"CA", X"D0", X"F7", X"CA", 
        X"9A", X"20", X"71", X"F0", X"D8", X"A9", X"00", X"85", 
        X"5B", X"20", X"CE", X"F0", X"A2", X"0F", X"86", X"58", 
        X"86", X"59", X"20", X"E5", X"FE", X"A9", X"3F", X"20", 
        X"EF", X"FF", X"20", X"E0", X"FE", X"20", X"EA", X"FE", 
        X"C9", X"08", X"F0", X"E0", X"C9", X"0D", X"F0", X"08", 
        X"20", X"EF", X"FF", X"95", X"00", X"E8", X"D0", X"ED", 
        X"A5", X"0F", X"F0", X"D0", X"A5", X"10", X"F0", X"04", 
        X"C9", X"20", X"D0", X"0C", X"A2", X"0D", X"BD", X"27", 
        X"FD", X"C5", X"0F", X"F0", X"0E", X"CA", X"D0", X"F6", 
        X"48", X"48", X"A0", X"03", X"68", X"68", X"20", X"69", 
        X"F4", X"D0", X"B1", X"20", X"D6", X"F0", X"4C", X"1C", 
        X"F0", X"A9", X"00", X"A8", X"85", X"FE", X"91", X"FE", 
        X"A5", X"FF", X"85", X"FD", X"A9", X"00", X"85", X"FA", 
        X"85", X"FB", X"85", X"FC", X"60", X"20", X"71", X"F0", 
        X"A5", X"11", X"D0", X"02", X"A9", X"01", X"91", X"FE", 
        X"60", X"20", X"AB", X"F0", X"F0", X"CC", X"20", X"E5", 
        X"FE", X"A5", X"3F", X"A6", X"3E", X"4C", X"67", X"FB", 
        X"20", X"AB", X"F0", X"F0", X"BD", X"20", X"E5", X"FE", 
        X"6C", X"3E", X"00", X"A2", X"02", X"B5", X"0F", X"F0", 
        X"08", X"48", X"20", X"D3", X"F7", X"68", X"E8", X"F0", 
        X"AB", X"60", X"A5", X"F5", X"85", X"3E", X"A5", X"F6", 
        X"85", X"3F", X"60", X"A5", X"3E", X"85", X"F5", X"A5", 
        X"3F", X"85", X"F6", X"60", X"A9", X"20", X"A2", X"27", 
        X"95", X"FF", X"CA", X"D0", X"FB", X"60", X"BD", X"34", 
        X"FD", X"48", X"BD", X"41", X"FD", X"48", X"60", X"20", 
        X"71", X"F0", X"4C", X"58", X"F1", X"20", X"78", X"F0", 
        X"20", X"1D", X"F1", X"F0", X"03", X"20", X"53", X"F2", 
        X"A0", X"00", X"B1", X"FC", X"F0", X"0E", X"20", X"72", 
        X"F2", X"20", X"DC", X"F4", X"AD", X"11", X"D0", X"10", 
        X"EF", X"AD", X"10", X"D0", X"60", X"20", X"4F", X"F2", 
        X"20", X"E5", X"FE", X"A2", X"04", X"B5", X"FB", X"20", 
        X"DC", X"FF", X"E0", X"03", X"D0", X"03", X"20", X"B9", 
        X"FE", X"CA", X"D0", X"F1", X"60", X"A0", X"00", X"84", 
        X"30", X"A2", X"01", X"B5", X"0F", X"F0", X"25", X"C9", 
        X"20", X"F0", X"07", X"C9", X"24", X"F0", X"03", X"E8", 
        X"D0", X"F1", X"E6", X"30", X"A9", X"24", X"95", X"0F", 
        X"20", X"5B", X"F9", X"E8", X"F0", X"5F", X"A5", X"3E", 
        X"99", X"54", X"00", X"C8", X"A5", X"3F", X"99", X"54", 
        X"00", X"C8", X"D0", X"D7", X"A4", X"30", X"60", X"20", 
        X"1D", X"F1", X"88", X"D0", X"48", X"20", X"C7", X"F1", 
        X"20", X"1D", X"F1", X"E8", X"F0", X"3F", X"98", X"D0", 
        X"06", X"20", X"4F", X"F2", X"18", X"90", X"03", X"20", 
        X"53", X"F2", X"20", X"DE", X"F2", X"E0", X"FF", X"F0", 
        X"AB", X"86", X"2F", X"A5", X"FD", X"85", X"51", X"85", 
        X"53", X"A5", X"FC", X"85", X"50", X"18", X"65", X"2F", 
        X"85", X"52", X"90", X"02", X"E6", X"53", X"20", X"A0", 
        X"F1", X"20", X"25", X"F2", X"A0", X"00", X"B9", X"00", 
        X"00", X"91", X"FC", X"C8", X"C4", X"2F", X"D0", X"F6", 
        X"20", X"DC", X"F4", X"D0", X"CD", X"4C", X"62", X"F0", 
        X"A2", X"FC", X"B5", X"FE", X"48", X"E8", X"D0", X"FA", 
        X"20", X"4F", X"F2", X"38", X"A5", X"FC", X"E5", X"50", 
        X"85", X"54", X"A5", X"FD", X"E5", X"51", X"85", X"55", 
        X"E6", X"54", X"D0", X"02", X"E6", X"55", X"A2", X"04", 
        X"68", X"95", X"F9", X"CA", X"D0", X"FA", X"60", X"20", 
        X"1D", X"F1", X"F0", X"D1", X"84", X"30", X"20", X"53", 
        X"F2", X"E0", X"FF", X"F0", X"C8", X"A5", X"FC", X"85", 
        X"52", X"A5", X"FD", X"85", X"53", X"A5", X"30", X"4A", 
        X"F0", X"0C", X"A6", X"57", X"A4", X"56", X"E4", X"55", 
        X"D0", X"02", X"C4", X"54", X"90", X"AF", X"C8", X"D0", 
        X"01", X"E8", X"86", X"55", X"84", X"54", X"20", X"53", 
        X"F2", X"A5", X"FC", X"85", X"50", X"A5", X"FD", X"85", 
        X"51", X"20", X"A0", X"F1", X"A0", X"00", X"A6", X"55", 
        X"F0", X"0E", X"B1", X"50", X"91", X"52", X"C8", X"D0", 
        X"F9", X"E6", X"51", X"E6", X"53", X"CA", X"D0", X"F2", 
        X"A6", X"54", X"F0", X"08", X"B1", X"50", X"91", X"52", 
        X"C8", X"CA", X"D0", X"F8", X"60", X"A6", X"55", X"18", 
        X"8A", X"65", X"51", X"85", X"51", X"18", X"8A", X"65", 
        X"53", X"85", X"53", X"E8", X"A4", X"54", X"F0", X"0E", 
        X"88", X"F0", X"07", X"B1", X"50", X"91", X"52", X"88", 
        X"D0", X"F9", X"B1", X"50", X"91", X"52", X"88", X"C6", 
        X"51", X"C6", X"53", X"CA", X"D0", X"ED", X"60", X"A9", 
        X"FF", X"85", X"55", X"20", X"78", X"F0", X"A4", X"54", 
        X"C4", X"FA", X"D0", X"06", X"A6", X"55", X"E4", X"FB", 
        X"F0", X"51", X"A0", X"FF", X"C8", X"B1", X"FC", X"D0", 
        X"FB", X"98", X"F0", X"45", X"C8", X"20", X"DC", X"F4", 
        X"D0", X"E4", X"20", X"E5", X"FE", X"86", X"2F", X"20", 
        X"EE", X"F3", X"C8", X"20", X"D6", X"FE", X"A2", X"00", 
        X"B5", X"04", X"F0", X"06", X"20", X"EF", X"FF", X"E8", 
        X"D0", X"F6", X"A6", X"2F", X"60", X"20", X"EA", X"FE", 
        X"C9", X"09", X"D0", X"02", X"A9", X"20", X"C9", X"20", 
        X"10", X"1A", X"A8", X"68", X"68", X"68", X"68", X"C0", 
        X"08", X"F0", X"3B", X"C0", X"0D", X"D0", X"0A", X"E0", 
        X"04", X"F0", X"29", X"A9", X"00", X"95", X"00", X"F0", 
        X"5C", X"A2", X"FF", X"60", X"E0", X"27", X"10", X"1A", 
        X"C9", X"5E", X"10", X"16", X"38", X"60", X"C9", X"2E", 
        X"F0", X"FA", X"C9", X"30", X"30", X"0C", X"C9", X"3A", 
        X"30", X"F2", X"C9", X"41", X"30", X"04", X"C9", X"5B", 
        X"30", X"EA", X"18", X"60", X"A9", X"02", X"AA", X"85", 
        X"00", X"A9", X"00", X"85", X"01", X"60", X"20", X"CC", 
        X"F0", X"A9", X"00", X"85", X"1D", X"20", X"E5", X"FE", 
        X"20", X"D6", X"FE", X"A2", X"04", X"A9", X"0A", X"20", 
        X"9C", X"F3", X"20", X"C4", X"F3", X"A5", X"04", X"C9", 
        X"3B", X"F0", X"0D", X"A9", X"0E", X"20", X"9C", X"F3", 
        X"20", X"C4", X"F3", X"A9", X"1D", X"20", X"9C", X"F3", 
        X"A9", X"00", X"20", X"9C", X"F3", X"A2", X"00", X"86", 
        X"51", X"A9", X"20", X"85", X"55", X"A9", X"04", X"85", 
        X"50", X"A9", X"01", X"85", X"54", X"20", X"D7", X"F3", 
        X"A4", X"04", X"C0", X"3B", X"D0", X"04", X"A9", X"0B", 
        X"D0", X"5F", X"8A", X"48", X"18", X"66", X"56", X"A2", 
        X"03", X"38", X"B5", X"0A", X"E9", X"40", X"A0", X"05", 
        X"4A", X"66", X"56", X"66", X"57", X"88", X"D0", X"F8", 
        X"CA", X"D0", X"EE", X"A2", X"38", X"BD", X"E8", X"FB", 
        X"C5", X"56", X"D0", X"07", X"BD", X"20", X"FC", X"C5", 
        X"57", X"F0", X"03", X"CA", X"D0", X"EF", X"CA", X"8A", 
        X"C9", X"FF", X"D0", X"19", X"A5", X"0B", X"C9", X"2E", 
        X"D0", X"0C", X"A2", X"05", X"A5", X"0C", X"DD", X"4E", 
        X"FD", X"F0", X"09", X"CA", X"D0", X"F8", X"68", X"A0", 
        X"01", X"4C", X"69", X"F4", X"CA", X"A8", X"C8", X"68", 
        X"AA", X"94", X"00", X"E8", X"A9", X"0F", X"85", X"50", 
        X"20", X"D7", X"F3", X"86", X"2F", X"E6", X"2F", X"A9", 
        X"1D", X"85", X"50", X"A9", X"00", X"85", X"54", X"85", 
        X"55", X"20", X"D7", X"F3", X"E4", X"2F", X"D0", X"03", 
        X"CA", X"95", X"FF", X"60", X"85", X"54", X"20", X"8D", 
        X"F2", X"90", X"FB", X"20", X"EF", X"FF", X"95", X"00", 
        X"E8", X"C9", X"20", X"F0", X"05", X"E4", X"54", X"D0", 
        X"ED", X"60", X"A5", X"54", X"F0", X"E8", X"E4", X"54", 
        X"F0", X"F7", X"A9", X"20", X"95", X"00", X"20", X"EF", 
        X"FF", X"E8", X"D0", X"EE", X"B5", X"FF", X"C9", X"20", 
        X"F0", X"07", X"20", X"8D", X"F2", X"C9", X"20", X"D0", 
        X"F9", X"95", X"00", X"E8", X"4C", X"EF", X"FF", X"A0", 
        X"00", X"B1", X"50", X"F0", X"0B", X"C5", X"55", X"F0", 
        X"07", X"95", X"00", X"E8", X"E6", X"50", X"D0", X"F1", 
        X"A5", X"54", X"95", X"00", X"E8", X"60", X"20", X"CC", 
        X"F0", X"A0", X"00", X"A2", X"04", X"B1", X"FC", X"F0", 
        X"4D", X"C9", X"02", X"D0", X"05", X"C8", X"A9", X"00", 
        X"F0", X"46", X"C9", X"01", X"F0", X"06", X"95", X"00", 
        X"E8", X"C8", X"D0", X"E9", X"A5", X"04", X"C9", X"3B", 
        X"D0", X"04", X"A2", X"0B", X"D0", X"2D", X"C8", X"B1", 
        X"FC", X"AA", X"CA", X"86", X"3C", X"E0", X"38", X"10", 
        X"09", X"98", X"48", X"20", X"99", X"FA", X"68", X"A8", 
        X"D0", X"06", X"86", X"0C", X"A9", X"2E", X"85", X"0B", 
        X"C8", X"A2", X"0F", X"B1", X"FC", X"F0", X"11", X"C9", 
        X"01", X"D0", X"05", X"C8", X"A2", X"1D", X"D0", X"F3", 
        X"95", X"00", X"E8", X"C8", X"D0", X"ED", X"A2", X"FE", 
        X"95", X"00", X"60", X"20", X"94", X"F4", X"20", X"E5", 
        X"FE", X"20", X"F8", X"F5", X"20", X"B8", X"F4", X"E8", 
        X"F0", X"0F", X"E0", X"FF", X"D0", X"F6", X"E6", X"58", 
        X"20", X"10", X"F6", X"E8", X"F0", X"03", X"4C", X"F8", 
        X"F5", X"20", X"E5", X"FE", X"A2", X"05", X"BD", X"53", 
        X"FD", X"20", X"EF", X"FF", X"CA", X"D0", X"F7", X"98", 
        X"18", X"8A", X"69", X"03", X"88", X"D0", X"FB", X"A8", 
        X"A2", X"03", X"B9", X"56", X"FD", X"20", X"EF", X"FF", 
        X"C8", X"CA", X"D0", X"F6", X"CA", X"A5", X"59", X"D0", 
        X"26", X"4C", X"72", X"F2", X"20", X"78", X"F0", X"85", 
        X"58", X"85", X"EB", X"85", X"E9", X"85", X"F5", X"A5", 
        X"F8", X"85", X"F6", X"20", X"EB", X"F5", X"86", X"EA", 
        X"A9", X"00", X"85", X"2B", X"85", X"29", X"85", X"46", 
        X"A4", X"F9", X"C8", X"84", X"2A", X"84", X"47", X"60", 
        X"20", X"EE", X"F3", X"E0", X"FE", X"F0", X"1D", X"E0", 
        X"04", X"F0", X"18", X"A9", X"00", X"85", X"59", X"85", 
        X"58", X"85", X"5A", X"20", X"44", X"F5", X"E0", X"FF", 
        X"F0", X"1D", X"A0", X"00", X"B1", X"FC", X"F0", X"03", 
        X"C8", X"D0", X"F9", X"C8", X"A5", X"FC", X"84", X"44", 
        X"18", X"65", X"44", X"85", X"FC", X"90", X"02", X"E6", 
        X"FD", X"E6", X"FA", X"D0", X"02", X"E6", X"FB", X"60", 
        X"A4", X"3C", X"B9", X"73", X"FC", X"A6", X"3D", X"18", 
        X"7D", X"AB", X"FC", X"E0", X"0B", X"F0", X"0E", X"E0", 
        X"02", X"D0", X"11", X"C0", X"28", X"30", X"0D", X"C0", 
        X"30", X"B0", X"09", X"69", X"08", X"C0", X"35", X"D0", 
        X"03", X"18", X"69", X"04", X"20", X"2F", X"F5", X"C9", 
        X"00", X"D0", X"03", X"20", X"2F", X"F5", X"8A", X"F0", 
        X"CE", X"CA", X"F0", X"CB", X"A5", X"3E", X"E0", X"08", 
        X"30", X"05", X"20", X"2F", X"F5", X"A5", X"3F", X"A0", 
        X"00", X"91", X"F5", X"E6", X"F5", X"D0", X"02", X"E6", 
        X"F6", X"60", X"20", X"A9", X"F6", X"E0", X"FF", X"D0", 
        X"AF", X"A0", X"02", X"60", X"A5", X"04", X"C9", X"3B", 
        X"F0", X"A5", X"A6", X"0B", X"E0", X"2E", X"D0", X"0D", 
        X"A6", X"0C", X"E0", X"4D", X"D0", X"03", X"4C", X"B6", 
        X"F5", X"E0", X"3D", X"F0", X"47", X"C9", X"20", X"F0", 
        X"03", X"20", X"DF", X"F8", X"A5", X"0B", X"C9", X"2E", 
        X"D0", X"D0", X"A2", X"00", X"A5", X"0C", X"C9", X"53", 
        X"F0", X"19", X"85", X"58", X"20", X"7A", X"F7", X"E8", 
        X"F0", X"0C", X"A5", X"3E", X"A6", X"0C", X"E0", X"57", 
        X"F0", X"A8", X"A6", X"3F", X"F0", X"A9", X"A0", X"03", 
        X"A2", X"FF", X"60", X"B5", X"0F", X"C9", X"27", X"D0", 
        X"F5", X"E8", X"B5", X"0F", X"F0", X"F0", X"C9", X"27", 
        X"F0", X"09", X"20", X"2F", X"F5", X"E0", X"0E", X"D0", 
        X"F0", X"F0", X"E3", X"60", X"85", X"58", X"20", X"C2", 
        X"F2", X"90", X"DB", X"A2", X"00", X"20", X"7A", X"F7", 
        X"E8", X"F0", X"D3", X"4C", X"E2", X"F8", X"20", X"C2", 
        X"F2", X"90", X"CB", X"A0", X"00", X"A5", X"0F", X"F0", 
        X"14", X"C9", X"20", X"F0", X"10", X"20", X"F6", X"F5", 
        X"A2", X"00", X"A5", X"0F", X"20", X"5B", X"F9", X"E8", 
        X"F0", X"B4", X"20", X"C3", X"F0", X"20", X"DF", X"F8", 
        X"E0", X"FF", X"F0", X"C7", X"20", X"10", X"F6", X"E0", 
        X"FF", X"F0", X"C0", X"20", X"C4", X"FE", X"A9", X"00", 
        X"20", X"F6", X"F5", X"A2", X"00", X"86", X"EE", X"86", 
        X"EC", X"A6", X"F9", X"86", X"ED", X"60", X"85", X"58", 
        X"A5", X"F6", X"A6", X"F5", X"A4", X"58", X"F0", X"0D", 
        X"48", X"20", X"B9", X"FE", X"68", X"E0", X"00", X"D0", 
        X"03", X"38", X"E9", X"01", X"CA", X"4C", X"67", X"FB", 
        X"A6", X"2B", X"F0", X"72", X"86", X"59", X"86", X"45", 
        X"A5", X"F5", X"48", X"A5", X"F6", X"48", X"20", X"A8", 
        X"F4", X"A0", X"00", X"A5", X"58", X"85", X"48", X"84", 
        X"5A", X"B1", X"46", X"C9", X"2E", X"D0", X"02", X"85", 
        X"58", X"B1", X"46", X"99", X"1D", X"00", X"C8", X"C0", 
        X"06", X"D0", X"F6", X"B1", X"46", X"85", X"F5", X"C8", 
        X"B1", X"46", X"85", X"F6", X"C8", X"B1", X"46", X"85", 
        X"54", X"20", X"7E", X"F8", X"E0", X"FF", X"F0", X"47", 
        X"A5", X"5A", X"F0", X"04", X"A5", X"54", X"91", X"50", 
        X"20", X"C3", X"F7", X"A0", X"00", X"B1", X"F5", X"29", 
        X"1F", X"C9", X"10", X"F0", X"22", X"20", X"33", X"F5", 
        X"A5", X"3E", X"20", X"2A", X"F5", X"18", X"A5", X"46", 
        X"69", X"09", X"85", X"46", X"90", X"02", X"E6", X"47", 
        X"A5", X"48", X"85", X"58", X"C6", X"45", X"D0", X"A1", 
        X"68", X"85", X"F6", X"68", X"85", X"F5", X"60", X"20", 
        X"62", X"F7", X"E0", X"FF", X"F0", X"09", X"A0", X"01", 
        X"A5", X"3E", X"91", X"F5", X"4C", X"6D", X"F6", X"A0", 
        X"00", X"20", X"E0", X"FE", X"B1", X"46", X"20", X"EF", 
        X"FF", X"C8", X"C0", X"06", X"D0", X"F6", X"88", X"D0", 
        X"D7", X"A2", X"FF", X"86", X"3D", X"A5", X"3C", X"A6", 
        X"0F", X"F0", X"04", X"E0", X"20", X"D0", X"0E", X"A2", 
        X"00", X"20", X"3D", X"F7", X"E0", X"FF", X"D0", X"35", 
        X"A2", X"01", X"4C", X"3D", X"F7", X"E0", X"23", X"F0", 
        X"0E", X"A2", X"03", X"20", X"3D", X"F7", X"E0", X"FF", 
        X"F0", X"24", X"A5", X"0F", X"4C", X"4F", X"F7", X"C9", 
        X"2C", X"F0", X"71", X"A2", X"02", X"C9", X"35", X"F0", 
        X"07", X"20", X"3D", X"F7", X"E0", X"FF", X"F0", X"0D", 
        X"86", X"3D", X"CA", X"20", X"7A", X"F7", X"E8", X"F0", 
        X"5B", X"A5", X"3F", X"D0", X"57", X"60", X"A2", X"00", 
        X"A5", X"0F", X"C9", X"28", X"D0", X"01", X"E8", X"20", 
        X"D3", X"F7", X"E0", X"FF", X"F0", X"EF", X"20", X"9C", 
        X"F9", X"E0", X"FF", X"F0", X"E8", X"86", X"3D", X"E0", 
        X"06", X"D0", X"0E", X"A5", X"3C", X"C9", X"28", X"90", 
        X"08", X"C9", X"30", X"B0", X"04", X"A2", X"0B", X"D0", 
        X"28", X"A0", X"06", X"B9", X"15", X"FD", X"C5", X"3C", 
        X"D0", X"0E", X"BE", X"1B", X"FD", X"E4", X"3D", X"F0", 
        X"18", X"BE", X"21", X"FD", X"E4", X"3D", X"F0", X"11", 
        X"88", X"D0", X"E8", X"A6", X"3D", X"A5", X"3C", X"DD", 
        X"59", X"FC", X"90", X"08", X"DD", X"66", X"FC", X"B0", 
        X"03", X"86", X"3D", X"60", X"A2", X"FF", X"60", X"A2", 
        X"00", X"86", X"3E", X"86", X"3F", X"C9", X"2A", X"D0", 
        X"06", X"20", X"BA", X"F0", X"20", X"FD", X"F7", X"20", 
        X"D3", X"F7", X"38", X"A5", X"3E", X"E5", X"F5", X"85", 
        X"3E", X"A5", X"3F", X"E5", X"F6", X"85", X"3F", X"F0", 
        X"04", X"E6", X"3F", X"D0", X"D7", X"C6", X"3E", X"C6", 
        X"3E", X"60", X"B5", X"0F", X"F0", X"CE", X"C9", X"27", 
        X"F0", X"03", X"4C", X"D3", X"F7", X"E8", X"A9", X"00", 
        X"85", X"3F", X"B5", X"0F", X"85", X"3E", X"E8", X"B5", 
        X"0F", X"C9", X"27", X"D0", X"B7", X"E8", X"B5", X"0F", 
        X"F0", X"7C", X"C9", X"20", X"F0", X"78", X"48", X"E8", 
        X"B5", X"0F", X"20", X"51", X"FA", X"E0", X"FF", X"D0", 
        X"02", X"68", X"60", X"85", X"54", X"68", X"C9", X"2B", 
        X"F0", X"09", X"A5", X"54", X"18", X"49", X"FF", X"69", 
        X"01", X"85", X"54", X"A5", X"5A", X"F0", X"04", X"A5", 
        X"54", X"91", X"50", X"A5", X"54", X"10", X"02", X"C6", 
        X"3F", X"18", X"65", X"3E", X"85", X"3E", X"90", X"02", 
        X"E6", X"3F", X"60", X"86", X"56", X"B5", X"0F", X"C9", 
        X"3C", X"F0", X"04", X"C9", X"3E", X"D0", X"05", X"85", 
        X"58", X"E8", X"B5", X"0F", X"20", X"BE", X"F2", X"B0", 
        X"09", X"20", X"5B", X"F9", X"E0", X"FF", X"F0", X"24", 
        X"D0", X"0B", X"86", X"2F", X"20", X"60", X"F8", X"E0", 
        X"FF", X"F0", X"1B", X"A6", X"2F", X"E8", X"B5", X"0F", 
        X"20", X"BE", X"F2", X"B0", X"F8", X"C9", X"2B", X"F0", 
        X"04", X"C9", X"2D", X"D0", X"0A", X"20", X"9E", X"F7", 
        X"E0", X"FF", X"D0", X"E9", X"A0", X"03", X"60", X"A0", 
        X"00", X"A5", X"58", X"C9", X"3C", X"F0", X"08", X"C9", 
        X"3E", X"D0", X"06", X"A5", X"3F", X"85", X"3E", X"84", 
        X"3F", X"B5", X"0F", X"99", X"1D", X"00", X"F0", X"0A", 
        X"C9", X"20", X"F0", X"06", X"E8", X"C8", X"E0", X"0E", 
        X"D0", X"EF", X"A9", X"00", X"99", X"1D", X"00", X"A4", 
        X"56", X"A9", X"24", X"99", X"0F", X"00", X"C8", X"A5", 
        X"3F", X"F0", X"03", X"20", X"82", X"FA", X"A5", X"3E", 
        X"20", X"82", X"FA", X"A2", X"00", X"B5", X"1D", X"99", 
        X"0F", X"00", X"F0", X"BA", X"E8", X"C8", X"D0", X"F5", 
        X"A0", X"00", X"C0", X"06", X"F0", X"18", X"20", X"BE", 
        X"F2", X"90", X"09", X"99", X"1D", X"00", X"E8", X"B5", 
        X"0F", X"C8", X"D0", X"EE", X"A9", X"20", X"99", X"1D", 
        X"00", X"C8", X"C0", X"06", X"D0", X"F8", X"A9", X"1D", 
        X"85", X"42", X"A2", X"00", X"86", X"43", X"A9", X"06", 
        X"85", X"2E", X"A9", X"08", X"85", X"2D", X"A5", X"1D", 
        X"C9", X"2E", X"F0", X"11", X"20", X"8A", X"F9", X"F0", 
        X"13", X"A0", X"06", X"B1", X"40", X"85", X"3E", X"C8", 
        X"B1", X"40", X"85", X"3F", X"60", X"A2", X"03", X"20", 
        X"8A", X"F9", X"D0", X"ED", X"A5", X"58", X"D0", X"4F", 
        X"20", X"BA", X"F0", X"A5", X"2A", X"85", X"51", X"A5", 
        X"29", X"A6", X"2B", X"F0", X"0A", X"18", X"69", X"09", 
        X"90", X"02", X"E6", X"51", X"CA", X"D0", X"F6", X"85", 
        X"50", X"E6", X"2B", X"A5", X"2B", X"C9", X"55", X"10", 
        X"32", X"A9", X"1D", X"85", X"5A", X"85", X"52", X"20", 
        X"43", X"F9", X"C8", X"8A", X"91", X"50", X"60", X"20", 
        X"BA", X"F0", X"A9", X"04", X"85", X"52", X"85", X"42", 
        X"A2", X"00", X"86", X"43", X"A9", X"06", X"85", X"2E", 
        X"A5", X"04", X"C9", X"2E", X"D0", X"02", X"A2", X"03", 
        X"20", X"8A", X"F9", X"F0", X"0B", X"68", X"68", X"A0", 
        X"05", X"D0", X"02", X"A0", X"04", X"A2", X"FF", X"60", 
        X"A6", X"04", X"E0", X"2E", X"F0", X"17", X"38", X"A5", 
        X"E9", X"E9", X"08", X"B0", X"02", X"C6", X"EA", X"85", 
        X"E9", X"E6", X"EB", X"F0", X"E6", X"85", X"50", X"A5", 
        X"EA", X"85", X"51", X"D0", X"1E", X"A5", X"ED", X"85", 
        X"51", X"A5", X"EC", X"A6", X"EE", X"F0", X"0A", X"18", 
        X"69", X"08", X"90", X"02", X"E6", X"51", X"CA", X"D0", 
        X"F6", X"85", X"50", X"E6", X"EE", X"A5", X"EE", X"C9", 
        X"20", X"10", X"C0", X"A0", X"00", X"84", X"53", X"A2", 
        X"06", X"B1", X"52", X"91", X"50", X"C8", X"CA", X"D0", 
        X"F8", X"A5", X"3E", X"91", X"50", X"C8", X"A5", X"3F", 
        X"91", X"50", X"60", X"C9", X"24", X"D0", X"A6", X"84", 
        X"1E", X"20", X"18", X"FA", X"E0", X"FF", X"F0", X"9D", 
        X"85", X"1D", X"A0", X"00", X"84", X"3F", X"CA", X"CA", 
        X"B5", X"0F", X"C9", X"24", X"F0", X"06", X"20", X"51", 
        X"FA", X"38", X"B0", X"03", X"20", X"6D", X"FA", X"99", 
        X"3E", X"00", X"C8", X"C4", X"1D", X"D0", X"E7", X"A4", 
        X"1E", X"60", X"B5", X"E9", X"85", X"40", X"B5", X"EA", 
        X"85", X"41", X"B5", X"EB", X"85", X"2C", X"20", X"2C", 
        X"FA", X"E0", X"FF", X"60", X"A2", X"00", X"A9", X"04", 
        X"B4", X"0F", X"C0", X"28", X"D0", X"04", X"18", X"69", 
        X"03", X"E8", X"48", X"20", X"18", X"FA", X"A8", X"CA", 
        X"A5", X"3C", X"C9", X"21", X"F0", X"04", X"C9", X"23", 
        X"D0", X"01", X"C8", X"68", X"E8", X"F0", X"56", X"88", 
        X"F0", X"03", X"18", X"69", X"06", X"A8", X"B5", X"0F", 
        X"F0", X"04", X"C9", X"20", X"D0", X"14", X"A5", X"0F", 
        X"C9", X"28", X"F0", X"41", X"C0", X"0F", X"10", X"3D", 
        X"C0", X"07", X"F0", X"39", X"30", X"01", X"88", X"98", 
        X"AA", X"60", X"C9", X"29", X"D0", X"0B", X"A9", X"20", 
        X"85", X"0F", X"E8", X"B5", X"0F", X"C9", X"2C", X"D0", 
        X"D5", X"B5", X"0F", X"C9", X"2C", X"D0", X"1E", X"E8", 
        X"B5", X"0F", X"C9", X"58", X"F0", X"0D", X"C9", X"59", 
        X"D0", X"13", X"A5", X"0F", X"C9", X"28", X"F0", X"0D", 
        X"95", X"0D", X"C8", X"C8", X"B5", X"0D", X"C9", X"29", 
        X"F0", X"03", X"E8", X"D0", X"B1", X"A2", X"FF", X"60", 
        X"A0", X"00", X"E8", X"C8", X"20", X"6E", X"FA", X"C9", 
        X"FF", X"D0", X"F7", X"98", X"4A", X"F0", X"EE", X"C9", 
        X"03", X"B0", X"EA", X"60", X"A5", X"2C", X"F0", X"E5", 
        X"A2", X"00", X"A0", X"FF", X"C8", X"C4", X"2E", X"F0", 
        X"DE", X"B1", X"40", X"D1", X"42", X"F0", X"F5", X"E8", 
        X"E4", X"2C", X"F0", X"D1", X"A5", X"40", X"18", X"65", 
        X"2D", X"85", X"40", X"90", X"E5", X"E6", X"41", X"B0", 
        X"E1", X"20", X"6E", X"FA", X"C9", X"FF", X"F0", X"BD", 
        X"48", X"20", X"6D", X"FA", X"CA", X"C9", X"FF", X"D0", 
        X"02", X"68", X"60", X"85", X"44", X"68", X"0A", X"0A", 
        X"0A", X"0A", X"65", X"44", X"60", X"E8", X"B5", X"0F", 
        X"49", X"30", X"C9", X"0A", X"90", X"08", X"69", X"88", 
        X"C9", X"FA", X"90", X"03", X"29", X"0F", X"60", X"A9", 
        X"FF", X"60", X"48", X"20", X"D6", X"FB", X"20", X"8A", 
        X"FA", X"68", X"29", X"0F", X"09", X"30", X"C9", X"3A", 
        X"90", X"02", X"69", X"06", X"99", X"0F", X"00", X"C8", 
        X"60", X"BD", X"E9", X"FB", X"85", X"56", X"BD", X"21", 
        X"FC", X"85", X"57", X"A2", X"00", X"A9", X"00", X"A0", 
        X"05", X"06", X"57", X"26", X"56", X"2A", X"88", X"D0", 
        X"F8", X"69", X"40", X"95", X"0B", X"A4", X"5B", X"F0", 
        X"03", X"20", X"EF", X"FF", X"E8", X"E0", X"03", X"D0", 
        X"E4", X"60", X"20", X"AB", X"F0", X"F0", X"03", X"20", 
        X"C3", X"F0", X"20", X"DC", X"FA", X"20", X"81", X"FB", 
        X"85", X"F5", X"84", X"F6", X"AD", X"11", X"D0", X"10", 
        X"F1", X"AD", X"10", X"D0", X"20", X"6E", X"FB", X"A1", 
        X"F5", X"A8", X"4A", X"90", X"09", X"6A", X"B0", X"14", 
        X"C9", X"A2", X"F0", X"10", X"29", X"87", X"4A", X"AA", 
        X"BD", X"B8", X"FC", X"90", X"03", X"20", X"D6", X"FB", 
        X"29", X"0F", X"D0", X"04", X"A0", X"80", X"A9", X"00", 
        X"AA", X"BD", X"FC", X"FC", X"85", X"29", X"29", X"03", 
        X"85", X"2A", X"98", X"20", X"90", X"FB", X"A0", X"00", 
        X"48", X"B1", X"F5", X"20", X"DC", X"FF", X"A2", X"01", 
        X"20", X"7A", X"FB", X"C4", X"2A", X"C8", X"90", X"F1", 
        X"A2", X"03", X"86", X"5B", X"C0", X"04", X"90", X"F0", 
        X"68", X"AA", X"20", X"99", X"FA", X"20", X"78", X"FB", 
        X"A4", X"2A", X"A2", X"06", X"E0", X"03", X"F0", X"1E", 
        X"06", X"29", X"90", X"0E", X"BD", X"09", X"FD", X"20", 
        X"EF", X"FF", X"BD", X"0F", X"FD", X"F0", X"03", X"20", 
        X"EF", X"FF", X"CA", X"D0", X"E7", X"86", X"5B", X"60", 
        X"88", X"30", X"E5", X"20", X"DC", X"FF", X"A5", X"29", 
        X"C9", X"E8", X"B1", X"F5", X"90", X"F2", X"20", X"84", 
        X"FB", X"AA", X"E8", X"D0", X"01", X"C8", X"98", X"20", 
        X"DC", X"FF", X"8A", X"4C", X"DC", X"FF", X"20", X"E5", 
        X"FE", X"A5", X"F6", X"A6", X"F5", X"20", X"67", X"FB", 
        X"A2", X"03", X"20", X"E0", X"FE", X"CA", X"D0", X"FA", 
        X"60", X"38", X"A5", X"2A", X"A4", X"F6", X"AA", X"10", 
        X"01", X"88", X"65", X"F5", X"90", X"01", X"C8", X"60", 
        X"85", X"54", X"29", X"8F", X"C9", X"8A", X"F0", X"43", 
        X"0A", X"C9", X"10", X"F0", X"37", X"A5", X"54", X"0A", 
        X"69", X"80", X"2A", X"0A", X"29", X"1F", X"69", X"20", 
        X"48", X"A5", X"54", X"29", X"9F", X"F0", X"1B", X"0A", 
        X"C9", X"20", X"F0", X"10", X"29", X"06", X"D0", X"2F", 
        X"68", X"29", X"07", X"C9", X"03", X"10", X"02", X"69", 
        X"02", X"69", X"1F", X"60", X"68", X"29", X"07", X"69", 
        X"18", X"60", X"68", X"AA", X"BD", X"B0", X"FB", X"60", 
        X"16", X"21", X"17", X"18", X"A5", X"54", X"4A", X"4A", 
        X"4A", X"4A", X"60", X"20", X"D4", X"FB", X"C9", X"0E", 
        X"D0", X"02", X"69", X"FD", X"69", X"08", X"60", X"68", 
        X"60", X"82", X"1B", X"83", X"99", X"82", X"1B", X"83", 
        X"99", X"21", X"A6", X"A0", X"1B", X"4B", X"1B", X"4B", 
        X"99", X"A6", X"A6", X"A0", X"A4", X"21", X"73", X"14", 
        X"95", X"95", X"14", X"13", X"15", X"15", X"10", X"10", 
        X"13", X"11", X"54", X"12", X"53", X"9D", X"61", X"1C", 
        X"1C", X"7C", X"0B", X"2B", X"09", X"9D", X"61", X"1B", 
        X"98", X"0C", X"93", X"64", X"93", X"9D", X"61", X"21", 
        X"4B", X"20", X"06", X"20", X"46", X"02", X"12", X"02", 
        X"52", X"72", X"42", X"72", X"2C", X"B2", X"08", X"B0", 
        X"48", X"02", X"26", X"70", X"F0", X"70", X"E0", X"96", 
        X"12", X"26", X"18", X"52", X"86", X"A6", X"C6", X"E6", 
        X"8A", X"62", X"E4", X"68", X"60", X"32", X"32", X"32", 
        X"30", X"82", X"88", X"E4", X"06", X"02", X"02", X"60", 
        X"86", X"D8", X"D8", X"E4", X"E4", X"30", X"30", X"46", 
        X"86", X"00", X"30", X"25", X"19", X"24", X"28", X"34", 
        X"28", X"28", X"21", X"28", X"28", X"23", X"19", X"34", 
        X"30", X"21", X"38", X"34", X"36", X"30", X"30", X"38", 
        X"34", X"30", X"24", X"08", X"18", X"28", X"38", X"48", 
        X"58", X"68", X"78", X"88", X"98", X"A8", X"B8", X"C8", 
        X"D8", X"E8", X"F8", X"8A", X"9A", X"AA", X"BA", X"CA", 
        X"EA", X"00", X"40", X"60", X"10", X"30", X"50", X"70", 
        X"90", X"B0", X"D0", X"F0", X"14", X"20", X"40", X"80", 
        X"A0", X"C0", X"E0", X"01", X"21", X"41", X"61", X"81", 
        X"A1", X"C1", X"E1", X"02", X"22", X"42", X"62", X"82", 
        X"A2", X"C2", X"E2", X"00", X"08", X"00", X"00", X"04", 
        X"14", X"14", X"00", X"10", X"0C", X"1C", X"18", X"2C", 
        X"04", X"20", X"54", X"30", X"0D", X"80", X"04", X"90", 
        X"03", X"22", X"54", X"33", X"0D", X"80", X"04", X"90", 
        X"04", X"20", X"54", X"33", X"0D", X"80", X"04", X"90", 
        X"04", X"20", X"54", X"3B", X"0D", X"80", X"04", X"90", 
        X"00", X"22", X"44", X"33", X"0D", X"C8", X"44", X"00", 
        X"11", X"22", X"44", X"33", X"0D", X"C8", X"44", X"A9", 
        X"01", X"22", X"44", X"33", X"0D", X"80", X"04", X"90", 
        X"01", X"22", X"44", X"33", X"0D", X"80", X"04", X"90", 
        X"26", X"31", X"87", X"9A", X"00", X"21", X"81", X"82", 
        X"00", X"00", X"59", X"4D", X"91", X"92", X"86", X"4A", 
        X"85", X"9D", X"2C", X"29", X"2C", X"23", X"28", X"24", 
        X"59", X"00", X"58", X"24", X"24", X"00", X"22", X"24", 
        X"25", X"35", X"36", X"37", X"04", X"05", X"05", X"02", 
        X"05", X"05", X"04", X"05", X"0A", X"0B", X"0A", X"0A", 
        X"4E", X"4C", X"58", X"45", X"4D", X"52", X"44", X"49", 
        X"21", X"24", X"41", X"56", X"50", X"F0", X"F0", X"F1", 
        X"F1", X"F1", X"F0", X"FA", X"F1", X"FF", X"FF", X"F4", 
        X"F0", X"F0", X"DE", X"E4", X"C6", X"4E", X"04", X"9F", 
        X"C1", X"57", X"1A", X"0E", X"4A", X"90", X"84", X"42", 
        X"57", X"53", X"3D", X"4D", X"20", X"3A", X"52", X"52", 
        X"45", X"4D", X"4E", X"45", X"41", X"44", X"44", X"53", 
        X"59", X"4E", X"4F", X"56", X"46", X"53", X"59", X"4D", 
        X"4E", X"45", X"53", X"53", X"45", X"57", X"20", X"4E", 
        X"45", X"4B", X"20", X"59", X"42", X"20", X"33", X"2E", 
        X"31", X"20", X"52", X"45", X"44", X"41", X"53", X"55", 
        X"52", X"4B", X"0D", X"50", X"53", X"59", X"58", X"41", 
        X"4C", X"48", X"43", X"5A", X"49", X"44", X"42", X"00", 
        X"56", X"4E", X"20", X"E5", X"FE", X"20", X"B9", X"FE", 
        X"20", X"BE", X"FE", X"A0", X"07", X"D9", X"82", X"FD", 
        X"F0", X"5C", X"88", X"D0", X"F8", X"C9", X"52", X"D0", 
        X"06", X"20", X"9F", X"FE", X"6C", X"F5", X"00", X"C9", 
        X"54", X"D0", X"3A", X"A2", X"08", X"BD", X"96", X"FE", 
        X"95", X"E0", X"CA", X"D0", X"F8", X"A1", X"F5", X"F0", 
        X"5D", X"A4", X"2A", X"C9", X"20", X"F0", X"75", X"C9", 
        X"60", X"F0", X"63", X"C9", X"4C", X"F0", X"78", X"C9", 
        X"6C", X"F0", X"75", X"C9", X"40", X"F0", X"53", X"29", 
        X"1F", X"49", X"14", X"C9", X"04", X"F0", X"02", X"B1", 
        X"F5", X"99", X"E0", X"00", X"88", X"10", X"F8", X"20", 
        X"9F", X"FE", X"4C", X"E0", X"00", X"C9", X"21", X"D0", 
        X"06", X"20", X"1B", X"FF", X"4C", X"1E", X"FE", X"C9", 
        X"24", X"D0", X"97", X"4C", X"0F", X"FF", X"A2", X"FE", 
        X"20", X"BE", X"FE", X"95", X"11", X"E8", X"D0", X"F8", 
        X"20", X"51", X"FA", X"99", X"EF", X"00", X"A6", X"F1", 
        X"9A", X"4C", X"1E", X"FE", X"28", X"20", X"AA", X"FE", 
        X"68", X"85", X"F5", X"68", X"85", X"F6", X"BA", X"86", 
        X"F1", X"20", X"57", X"FE", X"20", X"DC", X"FA", X"4C", 
        X"92", X"FD", X"18", X"68", X"85", X"F0", X"68", X"85", 
        X"F5", X"68", X"85", X"F6", X"20", X"82", X"FB", X"84", 
        X"F6", X"18", X"90", X"14", X"18", X"20", X"82", X"FB", 
        X"AA", X"98", X"48", X"8A", X"48", X"A0", X"02", X"18", 
        X"B1", X"F5", X"AA", X"88", X"B1", X"F5", X"86", X"F6", 
        X"85", X"F5", X"B0", X"F3", X"4C", X"1E", X"FE", X"20", 
        X"E5", X"FE", X"A2", X"05", X"BD", X"82", X"FD", X"20", 
        X"EF", X"FF", X"20", X"B9", X"FE", X"B5", X"EF", X"20", 
        X"DC", X"FF", X"20", X"E0", X"FE", X"CA", X"D0", X"EC", 
        X"A5", X"F0", X"A2", X"08", X"0A", X"90", X"08", X"48", 
        X"BD", X"89", X"FD", X"20", X"EF", X"FF", X"68", X"CA", 
        X"D0", X"F2", X"60", X"18", X"A0", X"01", X"B1", X"F5", 
        X"20", X"84", X"FB", X"85", X"F5", X"98", X"38", X"B0", 
        X"A1", X"20", X"AA", X"FE", X"38", X"B0", X"9D", X"EA", 
        X"EA", X"4C", X"91", X"FE", X"4C", X"83", X"FE", X"A5", 
        X"F0", X"48", X"A5", X"F4", X"A6", X"F3", X"A4", X"F2", 
        X"28", X"60", X"85", X"F4", X"86", X"F3", X"84", X"F2", 
        X"08", X"68", X"85", X"F0", X"BA", X"86", X"F1", X"D8", 
        X"60", X"A9", X"2D", X"4C", X"EF", X"FF", X"20", X"EA", 
        X"FE", X"4C", X"EF", X"FF", X"20", X"E5", X"FE", X"A2", 
        X"00", X"B5", X"04", X"20", X"EF", X"FF", X"E8", X"E0", 
        X"06", X"D0", X"F6", X"20", X"E0", X"FE", X"A5", X"FB", 
        X"20", X"E5", X"FF", X"A5", X"FA", X"20", X"DC", X"FF", 
        X"A9", X"20", X"4C", X"EF", X"FF", X"A9", X"0D", X"4C", 
        X"EF", X"FF", X"AD", X"11", X"D0", X"10", X"FB", X"AD", 
        X"10", X"D0", X"29", X"7F", X"60", X"00", X"00", X"00", 
        X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
        X"D8", X"58", X"A0", X"7F", X"8C", X"12", X"D0", X"A9", 
        X"A7", X"8D", X"11", X"D0", X"8D", X"13", X"D0", X"A9", 
        X"5C", X"20", X"EF", X"FF", X"20", X"1B", X"FF", X"90", 
        X"F6", X"B0", X"F9", X"20", X"E5", X"FE", X"A0", X"01", 
        X"88", X"30", X"F8", X"20", X"BE", X"FE", X"99", X"00", 
        X"02", X"C9", X"0D", X"F0", X"0B", X"C9", X"5F", X"F0", 
        X"EF", X"C9", X"1B", X"F0", X"DA", X"C8", X"10", X"EB", 
        X"A0", X"FF", X"A9", X"00", X"AA", X"0A", X"85", X"2B", 
        X"C8", X"B9", X"00", X"02", X"C9", X"0D", X"D0", X"02", 
        X"38", X"60", X"09", X"80", X"C9", X"AE", X"90", X"F0", 
        X"F0", X"EC", X"C9", X"BA", X"F0", X"E7", X"C9", X"D2", 
        X"F0", X"3D", X"86", X"28", X"86", X"29", X"84", X"2A", 
        X"B9", X"00", X"02", X"49", X"30", X"C9", X"0A", X"90", 
        X"06", X"69", X"88", X"C9", X"FA", X"90", X"11", X"0A", 
        X"0A", X"0A", X"0A", X"A2", X"04", X"0A", X"26", X"28", 
        X"26", X"29", X"CA", X"D0", X"F8", X"C8", X"D0", X"E0", 
        X"C4", X"2A", X"D0", X"02", X"18", X"60", X"24", X"2B", 
        X"50", X"10", X"A5", X"28", X"81", X"26", X"E6", X"26", 
        X"D0", X"AF", X"E6", X"27", X"4C", X"41", X"FF", X"6C", 
        X"24", X"00", X"30", X"27", X"A2", X"02", X"B5", X"27", 
        X"95", X"25", X"95", X"23", X"CA", X"D0", X"F7", X"D0", 
        X"12", X"20", X"E5", X"FE", X"A5", X"25", X"20", X"DC", 
        X"FF", X"A5", X"24", X"20", X"DC", X"FF", X"A9", X"3A", 
        X"20", X"EF", X"FF", X"20", X"E0", X"FE", X"A1", X"24", 
        X"20", X"DC", X"FF", X"86", X"2B", X"A5", X"24", X"C5", 
        X"28", X"A5", X"25", X"E5", X"29", X"B0", X"C5", X"E6", 
        X"24", X"D0", X"02", X"E6", X"25", X"A5", X"24", X"29", 
        X"07", X"10", X"CC", X"00", X"48", X"4A", X"4A", X"4A", 
        X"4A", X"20", X"E5", X"FF", X"68", X"29", X"0F", X"09", 
        X"30", X"C9", X"3A", X"90", X"02", X"69", X"06", X"2C", 
        X"12", X"D0", X"30", X"FB", X"8D", X"12", X"D0", X"60", 
        X"00", X"00", X"00", X"0F", X"00", X"FF", X"00", X"01"
    );
    
begin
    process(clock)
    begin
        if rising_edge(clock) then
            if cs_n = '0' then
                data_out <= rom(to_integer(unsigned(address)));
            end if;
        end if;
    end process;

end rtl;
