-- ============================================================================
-- Replica1_CPU_6800.vhd
-- Derived from Replica1_CPU_Template.vhd
-- 
-- CPU: MC6809 (Motorola 6809 8-bit processor)
-- Dependencies: None (uses standard IEEE libraries only)
-- Note: This creates a "6800-based Replica 1" - different instruction set!
-- https://opencores.org/projects/system09
-- ============================================================================

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity CPU_6809 is
	port (
		-- Clock and Reset
		main_clk    : in  std_logic;        -- Main system clock
		reset_n     : in  std_logic;        -- Active low reset
		cpu_reset_n : in  std_logic;        -- Active low cpu reset
		E           : out std_logic;        -- Phase 2 clock output (divided from main_clk)
		
		-- CPU Control Interface
		rw          : out std_logic;        -- Read/Write (1=Read, 0=Write)
		vma         : out std_logic;        -- Valid Memory Access
		sync        : out std_logic;        -- Instruction fetch cycle
		
		-- Address and Data Bus
		addr        : out std_logic_vector(15 downto 0);  -- Address bus
		data_in     : in  std_logic_vector(7 downto 0);   -- Data input
		data_out    : out std_logic_vector(7 downto 0);   -- Data output
		
		-- Interrupt Interface  
		nmi_n       : in  std_logic;        -- Non-maskable interrupt (active low)
		irq_n       : in  std_logic;        -- Interrupt request (active low)
		so_n        : in  std_logic := '1'; -- Set overflow (not used by 6800)
		
		-- wait states
		mrdy        : in  std_logic
	);
end CPU_6809;

architecture MC6809_impl of CPU_6809 is

	component cpu_clock_gen is
		 Port (
			  clk_4x  : in  STD_LOGIC;
			  reset_n : in  STD_LOGIC;
			  mrdy    : in  STD_LOGIC;       -- Memory Ready
			  clk_1x  : out STD_LOGIC;       -- CPU clock (stretched)
			  clk_2x  : out STD_LOGIC;       -- 2x clock for 6502 cores
			  stretch : out STD_LOGIC        -- '1' only when actually stretching
		 );
	end component;
	
	-- MC6809 Component (cpu09 core)
	component cpu09 is
		port (	
			clk      :	in std_logic;
			rst      :  in std_logic;
			vma      : out std_logic;
			addr     : out std_logic_vector(15 downto 0);
			rw       : out std_logic;
			data_out : out std_logic_vector(7 downto 0);
			data_in  :  in std_logic_vector(7 downto 0);
			irq      :  in std_logic;
			firq     :  in std_logic;
			nmi      :  in std_logic;
			halt     :  in std_logic;
			hold     :  in std_logic
			);
	end component;
	

	-- Internal signals
	signal data_bus      : std_logic_vector(7 downto 0);
	signal address_bus   : std_logic_vector(15 downto 0);
	signal cpu_data_out  : std_logic_vector(7 downto 0);

	-- MC6809 specific signals
	signal mc6809_rw     : std_logic;
	signal mc6809_vma    : std_logic;
	signal mc6809_clk    : std_logic;

begin


	clk: cpu_clock_gen port map(clk_4x  => main_clk,
						 			    reset_n => reset_n,
									    mrdy    => mrdy,
									    clk_1x  => mc6809_clk,
									    clk_2x  => open,
									    stretch => open);	
										 
										 
	E <= mc6809_clk;

	-- Input data bus assignment
	data_bus <= data_in;

	-- MC6809 Instantiation
	mc6800_inst: cpu09 
		port map(
			clk     => mc6809_clk,                 -- CPU09 uses 1x clock
			rst     => not cpu_reset_n,            -- MC6809 uses active high reset
			vma     => mc6809_vma,
			addr    => address_bus,
			rw      => mc6809_rw,
			data_out=> cpu_data_out,
			data_in => data_bus,
			irq     => not irq_n,                  -- MC6809 uses active high
			firq    => '0',                        -- no firq on apple 1
			nmi     => not nmi_n,                  -- MC6809 uses active high
			halt    => '0',                        -- No halt for Apple 1
			hold    => '0'                         -- No DMA for Apple 1
		);
		
	-- Note: 6809 VMA timing is different from 6502:
	-- - 6502: VMA = phi2 (address valid during phi2 high)
	-- - 6809: VMA is generated by CPU based on internal state

	-- Output assignments
	addr     <= address_bus;
	data_out <= cpu_data_out;
	rw       <= mc6809_rw;
	sync     <= '0';
	vma      <= mc6809_vma;

end MC6809_impl;